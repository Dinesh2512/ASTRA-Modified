module fir(
    input [31:0] inData,
    input clk,
    input reset,
    input sel,
    output [31:0] outData,
    output [111:0] pufout);

    wire VDD, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_6_, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, my_FIR_filter_firBlock_left_Y_in_0_, my_FIR_filter_firBlock_left_N257, my_FIR_filter_firBlock_left_N258, my_FIR_filter_firBlock_left_N259, my_FIR_filter_firBlock_left_N260, my_FIR_filter_firBlock_left_N261, my_FIR_filter_firBlock_left_N262, my_FIR_filter_firBlock_left_N263, my_FIR_filter_firBlock_left_N264, my_FIR_filter_firBlock_left_N265,
         my_FIR_filter_firBlock_left_N266, my_FIR_filter_firBlock_left_N267, my_FIR_filter_firBlock_left_N268, my_FIR_filter_firBlock_left_N269, my_FIR_filter_firBlock_left_N270, my_FIR_filter_firBlock_left_N271, my_FIR_filter_firBlock_left_N272, my_FIR_filter_firBlock_left_N273, my_FIR_filter_firBlock_left_N274, my_FIR_filter_firBlock_left_N275, my_FIR_filter_firBlock_left_N276,
         my_FIR_filter_firBlock_left_N277, my_FIR_filter_firBlock_left_N278, my_FIR_filter_firBlock_left_N279, my_FIR_filter_firBlock_left_N280, my_FIR_filter_firBlock_left_N281, my_FIR_filter_firBlock_left_N282, my_FIR_filter_firBlock_left_N283, my_FIR_filter_firBlock_left_N284, my_FIR_filter_firBlock_left_N285, my_FIR_filter_firBlock_left_N286, my_FIR_filter_firBlock_left_N287,
         my_FIR_filter_firBlock_left_N288, my_FIR_filter_firBlock_left_N225, my_FIR_filter_firBlock_left_N226, my_FIR_filter_firBlock_left_N227, my_FIR_filter_firBlock_left_N228, my_FIR_filter_firBlock_left_N229, my_FIR_filter_firBlock_left_N230, my_FIR_filter_firBlock_left_N231, my_FIR_filter_firBlock_left_N232, my_FIR_filter_firBlock_left_N233, my_FIR_filter_firBlock_left_N234,
         my_FIR_filter_firBlock_left_N235, my_FIR_filter_firBlock_left_N236, my_FIR_filter_firBlock_left_N237, my_FIR_filter_firBlock_left_N238, my_FIR_filter_firBlock_left_N239, my_FIR_filter_firBlock_left_N240, my_FIR_filter_firBlock_left_N241, my_FIR_filter_firBlock_left_N242, my_FIR_filter_firBlock_left_N243, my_FIR_filter_firBlock_left_N244, my_FIR_filter_firBlock_left_N245,
         my_FIR_filter_firBlock_left_N246, my_FIR_filter_firBlock_left_N247, my_FIR_filter_firBlock_left_N248, my_FIR_filter_firBlock_left_N249, my_FIR_filter_firBlock_left_N250, my_FIR_filter_firBlock_left_N251, my_FIR_filter_firBlock_left_N252, my_FIR_filter_firBlock_left_N253, my_FIR_filter_firBlock_left_N254, my_FIR_filter_firBlock_left_N255, my_FIR_filter_firBlock_left_N256,
         my_FIR_filter_firBlock_left_N193, my_FIR_filter_firBlock_left_N194, my_FIR_filter_firBlock_left_N195, my_FIR_filter_firBlock_left_N196, my_FIR_filter_firBlock_left_N197, my_FIR_filter_firBlock_left_N198, my_FIR_filter_firBlock_left_N199, my_FIR_filter_firBlock_left_N200, my_FIR_filter_firBlock_left_N201, my_FIR_filter_firBlock_left_N202, my_FIR_filter_firBlock_left_N203,
         my_FIR_filter_firBlock_left_N204, my_FIR_filter_firBlock_left_N205, my_FIR_filter_firBlock_left_N206, my_FIR_filter_firBlock_left_N207, my_FIR_filter_firBlock_left_N208, my_FIR_filter_firBlock_left_N209, my_FIR_filter_firBlock_left_N210, my_FIR_filter_firBlock_left_N211, my_FIR_filter_firBlock_left_N212, my_FIR_filter_firBlock_left_N213, my_FIR_filter_firBlock_left_N214,
         my_FIR_filter_firBlock_left_N215, my_FIR_filter_firBlock_left_N216, my_FIR_filter_firBlock_left_N217, my_FIR_filter_firBlock_left_N218, my_FIR_filter_firBlock_left_N219, my_FIR_filter_firBlock_left_N220, my_FIR_filter_firBlock_left_N221, my_FIR_filter_firBlock_left_N222, my_FIR_filter_firBlock_left_N223, my_FIR_filter_firBlock_left_N224, my_FIR_filter_firBlock_left_N161,
         my_FIR_filter_firBlock_left_N162, my_FIR_filter_firBlock_left_N163, my_FIR_filter_firBlock_left_N164, my_FIR_filter_firBlock_left_N165, my_FIR_filter_firBlock_left_N166, my_FIR_filter_firBlock_left_N167, my_FIR_filter_firBlock_left_N168, my_FIR_filter_firBlock_left_N169, my_FIR_filter_firBlock_left_N170, my_FIR_filter_firBlock_left_N171, my_FIR_filter_firBlock_left_N172,
         my_FIR_filter_firBlock_left_N173, my_FIR_filter_firBlock_left_N174, my_FIR_filter_firBlock_left_N175, my_FIR_filter_firBlock_left_N176, my_FIR_filter_firBlock_left_N177, my_FIR_filter_firBlock_left_N178, my_FIR_filter_firBlock_left_N179, my_FIR_filter_firBlock_left_N180, my_FIR_filter_firBlock_left_N181, my_FIR_filter_firBlock_left_N182, my_FIR_filter_firBlock_left_N183,
         my_FIR_filter_firBlock_left_N184, my_FIR_filter_firBlock_left_N185, my_FIR_filter_firBlock_left_N186, my_FIR_filter_firBlock_left_N187, my_FIR_filter_firBlock_left_N188, my_FIR_filter_firBlock_left_N189, my_FIR_filter_firBlock_left_N190, my_FIR_filter_firBlock_left_N191, my_FIR_filter_firBlock_left_N192, my_FIR_filter_firBlock_left_N129, my_FIR_filter_firBlock_left_N130,
         my_FIR_filter_firBlock_left_N131, my_FIR_filter_firBlock_left_N132, my_FIR_filter_firBlock_left_N133, my_FIR_filter_firBlock_left_N134, my_FIR_filter_firBlock_left_N135, my_FIR_filter_firBlock_left_N136, my_FIR_filter_firBlock_left_N137, my_FIR_filter_firBlock_left_N138, my_FIR_filter_firBlock_left_N139, my_FIR_filter_firBlock_left_N140, my_FIR_filter_firBlock_left_N141,
         my_FIR_filter_firBlock_left_N142, my_FIR_filter_firBlock_left_N143, my_FIR_filter_firBlock_left_N144, my_FIR_filter_firBlock_left_N145, my_FIR_filter_firBlock_left_N146, my_FIR_filter_firBlock_left_N147, my_FIR_filter_firBlock_left_N148, my_FIR_filter_firBlock_left_N149, my_FIR_filter_firBlock_left_N150, my_FIR_filter_firBlock_left_N151, my_FIR_filter_firBlock_left_N152,
         my_FIR_filter_firBlock_left_N153, my_FIR_filter_firBlock_left_N154, my_FIR_filter_firBlock_left_N155, my_FIR_filter_firBlock_left_N156, my_FIR_filter_firBlock_left_N157, my_FIR_filter_firBlock_left_N158, my_FIR_filter_firBlock_left_N159, my_FIR_filter_firBlock_left_N160, my_FIR_filter_firBlock_left_N97, my_FIR_filter_firBlock_left_N98, my_FIR_filter_firBlock_left_N99,
         my_FIR_filter_firBlock_left_N100, my_FIR_filter_firBlock_left_N101, my_FIR_filter_firBlock_left_N102, my_FIR_filter_firBlock_left_N103, my_FIR_filter_firBlock_left_N104, my_FIR_filter_firBlock_left_N105, my_FIR_filter_firBlock_left_N106, my_FIR_filter_firBlock_left_N107, my_FIR_filter_firBlock_left_N108, my_FIR_filter_firBlock_left_N109, my_FIR_filter_firBlock_left_N110,
         my_FIR_filter_firBlock_left_N111, my_FIR_filter_firBlock_left_N112, my_FIR_filter_firBlock_left_N113, my_FIR_filter_firBlock_left_N114, my_FIR_filter_firBlock_left_N115, my_FIR_filter_firBlock_left_N116, my_FIR_filter_firBlock_left_N117, my_FIR_filter_firBlock_left_N118, my_FIR_filter_firBlock_left_N119, my_FIR_filter_firBlock_left_N120, my_FIR_filter_firBlock_left_N121,
         my_FIR_filter_firBlock_left_N122, my_FIR_filter_firBlock_left_N123, my_FIR_filter_firBlock_left_N124, my_FIR_filter_firBlock_left_N125, my_FIR_filter_firBlock_left_N126, my_FIR_filter_firBlock_left_N127, my_FIR_filter_firBlock_left_N128, my_FIR_filter_firBlock_left_N65, my_FIR_filter_firBlock_left_N66, my_FIR_filter_firBlock_left_N67, my_FIR_filter_firBlock_left_N68,
         my_FIR_filter_firBlock_left_N69, my_FIR_filter_firBlock_left_N70, my_FIR_filter_firBlock_left_N71, my_FIR_filter_firBlock_left_N72, my_FIR_filter_firBlock_left_N73, my_FIR_filter_firBlock_left_N74, my_FIR_filter_firBlock_left_N75, my_FIR_filter_firBlock_left_N76, my_FIR_filter_firBlock_left_N77, my_FIR_filter_firBlock_left_N78, my_FIR_filter_firBlock_left_N79,
         my_FIR_filter_firBlock_left_N80, my_FIR_filter_firBlock_left_N81, my_FIR_filter_firBlock_left_N82, my_FIR_filter_firBlock_left_N83, my_FIR_filter_firBlock_left_N84, my_FIR_filter_firBlock_left_N85, my_FIR_filter_firBlock_left_N86, my_FIR_filter_firBlock_left_N87, my_FIR_filter_firBlock_left_N88, my_FIR_filter_firBlock_left_N89, my_FIR_filter_firBlock_left_N90,
         my_FIR_filter_firBlock_left_N91, my_FIR_filter_firBlock_left_N92, my_FIR_filter_firBlock_left_N93, my_FIR_filter_firBlock_left_N94, my_FIR_filter_firBlock_left_N95, my_FIR_filter_firBlock_left_N96, my_FIR_filter_firBlock_left_N33, my_FIR_filter_firBlock_left_N34, my_FIR_filter_firBlock_left_N35, my_FIR_filter_firBlock_left_N36, my_FIR_filter_firBlock_left_N37,
         my_FIR_filter_firBlock_left_N38, my_FIR_filter_firBlock_left_N39, my_FIR_filter_firBlock_left_N40, my_FIR_filter_firBlock_left_N41, my_FIR_filter_firBlock_left_N42, my_FIR_filter_firBlock_left_N43, my_FIR_filter_firBlock_left_N44, my_FIR_filter_firBlock_left_N45, my_FIR_filter_firBlock_left_N46, my_FIR_filter_firBlock_left_N47, my_FIR_filter_firBlock_left_N48,
         my_FIR_filter_firBlock_left_N49, my_FIR_filter_firBlock_left_N50, my_FIR_filter_firBlock_left_N51, my_FIR_filter_firBlock_left_N52, my_FIR_filter_firBlock_left_N53, my_FIR_filter_firBlock_left_N54, my_FIR_filter_firBlock_left_N55, my_FIR_filter_firBlock_left_N56, my_FIR_filter_firBlock_left_N57, my_FIR_filter_firBlock_left_N58, my_FIR_filter_firBlock_left_N59,
         my_FIR_filter_firBlock_left_N60, my_FIR_filter_firBlock_left_N61, my_FIR_filter_firBlock_left_N62, my_FIR_filter_firBlock_left_N63, my_FIR_filter_firBlock_left_N64, my_FIR_filter_firBlock_left_N1, my_FIR_filter_firBlock_left_N2, my_FIR_filter_firBlock_left_N3, my_FIR_filter_firBlock_left_N4, my_FIR_filter_firBlock_left_N5, my_FIR_filter_firBlock_left_N6,
         my_FIR_filter_firBlock_left_N7, my_FIR_filter_firBlock_left_N8, my_FIR_filter_firBlock_left_N9, my_FIR_filter_firBlock_left_N10, my_FIR_filter_firBlock_left_N11, my_FIR_filter_firBlock_left_N12, my_FIR_filter_firBlock_left_N13, my_FIR_filter_firBlock_left_N14, my_FIR_filter_firBlock_left_N15, my_FIR_filter_firBlock_left_N16, my_FIR_filter_firBlock_left_N17,
         my_FIR_filter_firBlock_left_N18, my_FIR_filter_firBlock_left_N19, my_FIR_filter_firBlock_left_N20, my_FIR_filter_firBlock_left_N21, my_FIR_filter_firBlock_left_N22, my_FIR_filter_firBlock_left_N23, my_FIR_filter_firBlock_left_N24, my_FIR_filter_firBlock_left_N25, my_FIR_filter_firBlock_left_N26, my_FIR_filter_firBlock_left_N27, my_FIR_filter_firBlock_left_N28,
         my_FIR_filter_firBlock_left_N29, my_FIR_filter_firBlock_left_N30, my_FIR_filter_firBlock_left_N31, my_FIR_filter_firBlock_left_N32, n317, n485, n483, n484, n482, n316, n315,
         n314, n313, n481, n480, n479, n478, n312, n311, n310, n309, n477,
         n476, n475, n474, n308, n307, n306, n305, n486, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_8_, n103, n571,
         n517, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_9_, n137, n570, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_10_, n473, n569, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_11_, n303, n568, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_12_,
         n138, n567, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_13_, n304, n566, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_14_, n565, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_15_, n564, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_16_, n563,
         my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_17_, n562, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_18_, n561, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_19_, n560, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_20_, n559, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_21_, n558, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_22_,
         n557, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_23_, n556, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_24_, n555, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_25_, n554, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_26_, n553, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_27_, n552,
         my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_28_, n551, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_29_, n550, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_30_, n549, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_31_, n548, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_32_, n547, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_33_,
         n546, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_34_, n545, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_35_, n544, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_36_, n543, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_37_, n542, my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_38_, n541,
         n298, n518, n276, n277, n278, n123, n124, n125, n126, n279, n280,
         n281, n282, n127, n128, n129, n130, n283, n284, n285, n286, n131,
         n132, n133, n134, n287, n288, n289, n290, n291, n292, n293, n467,
         n519, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n121, n122, n297, n520,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n466, n521, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n120, n296, n522, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n402, n465, n523, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n216, n295, n524, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n119, n464, n525, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n118, n186, n294, n516, n169, n170, n171, n105, n106, n107,
         n108, n172, n173, n174, n175, n109, n110, n111, n112, n176, n177,
         n178, n179, n113, n114, n115, n116, n180, n181, n182, n183, n184,
         n185, n117, n463, n104, n526, n344, n139, n343, n140, n342, n141,
         n341, n142, n340, n143, n339, n144, n338, n145, n337, n146, n336,
         n147, n335, n148, n334, n149, n333, n150, n332, n151, n331, n152,
         n330, n153, n329, n154, n328, n155, n327, n156, n326, n157, n325,
         n158, n324, n159, n323, n160, n322, n161, n321, n162, n320, n163,
         n460, n166, n462, n167, n461, n168, n319, n164, n318, n165, n136,
         n472, n302, n471, n301, n470, n300, n469, n135, n468, n299, n66,
         n572, n573, n99, n530, n100, n531, n101, n539, n540, n538, n102,
         n527, n575, n514, n487, n603, n515, n488, n602, n489, n601, n490,
         n600, n491, n599, n492, n598, n493, n597, n494, n596, n495, n595,
         n496, n594, n497, n593, n498, n592, n499, n591, n500, n590, n501,
         n589, n502, n588, n503, n587, n504, n586, n505, n585, n506, n584,
         n507, n583, n508, n582, n509, n581, n510, n580, n511, n579, n512,
         n578, n513, n577, n576, n604, n605, n574, n528, n529, n532, n533,
         n534, n535, n536, n537, puf_0_wire_0, puf_0_wire_1, puf_0_wire_2, puf_0_wire_5, puf_0_wire_6, puf_0_wire_7, puf_0_wire_8,
         puf_1_wire_0, puf_1_wire_1, puf_1_wire_2, puf_1_wire_5, puf_1_wire_6, puf_1_wire_7, puf_1_wire_8, puf_2_wire_0, puf_2_wire_1, puf_2_wire_2, puf_2_wire_5,
         puf_2_wire_6, puf_2_wire_7, puf_2_wire_8, puf_3_wire_0, puf_3_wire_1, puf_3_wire_2, puf_3_wire_5, puf_3_wire_6, puf_3_wire_7, puf_3_wire_8, puf_4_wire_0,
         puf_4_wire_1, puf_4_wire_2, puf_4_wire_5, puf_4_wire_6, puf_4_wire_7, puf_4_wire_8, puf_5_wire_0, puf_5_wire_1, puf_5_wire_2, puf_5_wire_5, puf_5_wire_6,
         puf_5_wire_7, puf_5_wire_8, puf_6_wire_0, puf_6_wire_1, puf_6_wire_2, puf_6_wire_5, puf_6_wire_6, puf_6_wire_7, puf_6_wire_8, puf_7_wire_0, puf_7_wire_1,
         puf_7_wire_2, puf_7_wire_5, puf_7_wire_6, puf_7_wire_7, puf_7_wire_8, puf_8_wire_0, puf_8_wire_1, puf_8_wire_2, puf_8_wire_5, puf_8_wire_6, puf_8_wire_7,
         puf_8_wire_8, puf_9_wire_0, puf_9_wire_1, puf_9_wire_2, puf_9_wire_5, puf_9_wire_6, puf_9_wire_7, puf_9_wire_8, puf_10_wire_0, puf_10_wire_1, puf_10_wire_2,
         puf_10_wire_5, puf_10_wire_6, puf_10_wire_7, puf_10_wire_8, puf_11_wire_0, puf_11_wire_1, puf_11_wire_2, puf_11_wire_5, puf_11_wire_6, puf_11_wire_7, puf_11_wire_8,
         puf_12_wire_0, puf_12_wire_1, puf_12_wire_2, puf_12_wire_5, puf_12_wire_6, puf_12_wire_7, puf_12_wire_8, puf_13_wire_0, puf_13_wire_1, puf_13_wire_2, puf_13_wire_5,
         puf_13_wire_6, puf_13_wire_7, puf_13_wire_8, puf_14_wire_0, puf_14_wire_1, puf_14_wire_2, puf_14_wire_5, puf_14_wire_6, puf_14_wire_7, puf_14_wire_8, puf_15_wire_0,
         puf_15_wire_1, puf_15_wire_2, puf_15_wire_5, puf_15_wire_6, puf_15_wire_7, puf_15_wire_8, puf_16_wire_0, puf_16_wire_1, puf_16_wire_2, puf_16_wire_5, puf_16_wire_6,
         puf_16_wire_7, puf_16_wire_8, puf_17_wire_0, puf_17_wire_1, puf_17_wire_2, puf_17_wire_5, puf_17_wire_6, puf_17_wire_7, puf_17_wire_8, puf_18_wire_0, puf_18_wire_1,
         puf_18_wire_2, puf_18_wire_5, puf_18_wire_6, puf_18_wire_7, puf_18_wire_8, puf_19_wire_0, puf_19_wire_1, puf_19_wire_2, puf_19_wire_5, puf_19_wire_6, puf_19_wire_7,
         puf_19_wire_8, puf_20_wire_0, puf_20_wire_1, puf_20_wire_2, puf_20_wire_5, puf_20_wire_6, puf_20_wire_7, puf_20_wire_8, puf_21_wire_0, puf_21_wire_1, puf_21_wire_2,
         puf_21_wire_5, puf_21_wire_6, puf_21_wire_7, puf_21_wire_8, puf_22_wire_0, puf_22_wire_1, puf_22_wire_2, puf_22_wire_5, puf_22_wire_6, puf_22_wire_7, puf_22_wire_8,
         puf_23_wire_0, puf_23_wire_1, puf_23_wire_2, puf_23_wire_5, puf_23_wire_6, puf_23_wire_7, puf_23_wire_8, puf_24_wire_0, puf_24_wire_1, puf_24_wire_2, puf_24_wire_5,
         puf_24_wire_6, puf_24_wire_7, puf_24_wire_8, puf_25_wire_0, puf_25_wire_1, puf_25_wire_2, puf_25_wire_5, puf_25_wire_6, puf_25_wire_7, puf_25_wire_8, puf_26_wire_0,
         puf_26_wire_1, puf_26_wire_2, puf_26_wire_5, puf_26_wire_6, puf_26_wire_7, puf_26_wire_8, puf_27_wire_0, puf_27_wire_1, puf_27_wire_2, puf_27_wire_5, puf_27_wire_6,
         puf_27_wire_7, puf_27_wire_8, puf_28_wire_0, puf_28_wire_1, puf_28_wire_2, puf_28_wire_5, puf_28_wire_6, puf_28_wire_7, puf_28_wire_8, puf_29_wire_0, puf_29_wire_1,
         puf_29_wire_2, puf_29_wire_5, puf_29_wire_6, puf_29_wire_7, puf_29_wire_8, puf_30_wire_0, puf_30_wire_1, puf_30_wire_2, puf_30_wire_5, puf_30_wire_6, puf_30_wire_7,
         puf_30_wire_8, puf_31_wire_0, puf_31_wire_1, puf_31_wire_2, puf_31_wire_5, puf_31_wire_6, puf_31_wire_7, puf_31_wire_8, puf_32_wire_0, puf_32_wire_1, puf_32_wire_2,
         puf_32_wire_5, puf_32_wire_6, puf_32_wire_7, puf_32_wire_8, puf_33_wire_0, puf_33_wire_1, puf_33_wire_2, puf_33_wire_5, puf_33_wire_6, puf_33_wire_7, puf_33_wire_8,
         puf_34_wire_0, puf_34_wire_1, puf_34_wire_2, puf_34_wire_5, puf_34_wire_6, puf_34_wire_7, puf_34_wire_8, puf_35_wire_0, puf_35_wire_1, puf_35_wire_2, puf_35_wire_5,
         puf_35_wire_6, puf_35_wire_7, puf_35_wire_8, puf_36_wire_0, puf_36_wire_1, puf_36_wire_2, puf_36_wire_5, puf_36_wire_6, puf_36_wire_7, puf_36_wire_8, puf_37_wire_0,
         puf_37_wire_1, puf_37_wire_2, puf_37_wire_5, puf_37_wire_6, puf_37_wire_7, puf_37_wire_8, puf_38_wire_0, puf_38_wire_1, puf_38_wire_2, puf_38_wire_5, puf_38_wire_6,
         puf_38_wire_7, puf_38_wire_8, puf_39_wire_0, puf_39_wire_1, puf_39_wire_2, puf_39_wire_5, puf_39_wire_6, puf_39_wire_7, puf_39_wire_8, puf_40_wire_0, puf_40_wire_1,
         puf_40_wire_2, puf_40_wire_5, puf_40_wire_6, puf_40_wire_7, puf_40_wire_8, puf_41_wire_0, puf_41_wire_1, puf_41_wire_2, puf_41_wire_5, puf_41_wire_6, puf_41_wire_7,
         puf_41_wire_8, puf_42_wire_0, puf_42_wire_1, puf_42_wire_2, puf_42_wire_5, puf_42_wire_6, puf_42_wire_7, puf_42_wire_8, puf_43_wire_0, puf_43_wire_1, puf_43_wire_2,
         puf_43_wire_5, puf_43_wire_6, puf_43_wire_7, puf_43_wire_8, puf_44_wire_0, puf_44_wire_1, puf_44_wire_2, puf_44_wire_5, puf_44_wire_6, puf_44_wire_7, puf_44_wire_8,
         puf_45_wire_0, puf_45_wire_1, puf_45_wire_2, puf_45_wire_5, puf_45_wire_6, puf_45_wire_7, puf_45_wire_8, puf_46_wire_0, puf_46_wire_1, puf_46_wire_2, puf_46_wire_5,
         puf_46_wire_6, puf_46_wire_7, puf_46_wire_8, puf_47_wire_0, puf_47_wire_1, puf_47_wire_2, puf_47_wire_5, puf_47_wire_6, puf_47_wire_7, puf_47_wire_8, puf_48_wire_0,
         puf_48_wire_1, puf_48_wire_2, puf_48_wire_5, puf_48_wire_6, puf_48_wire_7, puf_48_wire_8, puf_49_wire_0, puf_49_wire_1, puf_49_wire_2, puf_49_wire_5, puf_49_wire_6,
         puf_49_wire_7, puf_49_wire_8, puf_50_wire_0, puf_50_wire_1, puf_50_wire_2, puf_50_wire_5, puf_50_wire_6, puf_50_wire_7, puf_50_wire_8, puf_51_wire_0, puf_51_wire_1,
         puf_51_wire_2, puf_51_wire_5, puf_51_wire_6, puf_51_wire_7, puf_51_wire_8, puf_52_wire_0, puf_52_wire_1, puf_52_wire_2, puf_52_wire_5, puf_52_wire_6, puf_52_wire_7,
         puf_52_wire_8, puf_53_wire_0, puf_53_wire_1, puf_53_wire_2, puf_53_wire_5, puf_53_wire_6, puf_53_wire_7, puf_53_wire_8, puf_54_wire_0, puf_54_wire_1, puf_54_wire_2,
         puf_54_wire_5, puf_54_wire_6, puf_54_wire_7, puf_54_wire_8, puf_55_wire_0, puf_55_wire_1, puf_55_wire_2, puf_55_wire_5, puf_55_wire_6, puf_55_wire_7, puf_55_wire_8,
         puf_56_wire_0, puf_56_wire_1, puf_56_wire_2, puf_56_wire_5, puf_56_wire_6, puf_56_wire_7, puf_56_wire_8, puf_57_wire_0, puf_57_wire_1, puf_57_wire_2, puf_57_wire_5,
         puf_57_wire_6, puf_57_wire_7, puf_57_wire_8, puf_58_wire_0, puf_58_wire_1, puf_58_wire_2, puf_58_wire_5, puf_58_wire_6, puf_58_wire_7, puf_58_wire_8, puf_59_wire_0,
         puf_59_wire_1, puf_59_wire_2, puf_59_wire_5, puf_59_wire_6, puf_59_wire_7, puf_59_wire_8, puf_60_wire_0, puf_60_wire_1, puf_60_wire_2, puf_60_wire_5, puf_60_wire_6,
         puf_60_wire_7, puf_60_wire_8, puf_61_wire_0, puf_61_wire_1, puf_61_wire_2, puf_61_wire_5, puf_61_wire_6, puf_61_wire_7, puf_61_wire_8, puf_62_wire_0, puf_62_wire_1,
         puf_62_wire_2, puf_62_wire_5, puf_62_wire_6, puf_62_wire_7, puf_62_wire_8, puf_63_wire_0, puf_63_wire_1, puf_63_wire_2, puf_63_wire_5, puf_63_wire_6, puf_63_wire_7,
         puf_63_wire_8, puf_64_wire_0, puf_64_wire_1, puf_64_wire_2, puf_64_wire_5, puf_64_wire_6, puf_64_wire_7, puf_64_wire_8, puf_65_wire_0, puf_65_wire_1, puf_65_wire_2,
         puf_65_wire_5, puf_65_wire_6, puf_65_wire_7, puf_65_wire_8, puf_66_wire_0, puf_66_wire_1, puf_66_wire_2, puf_66_wire_5, puf_66_wire_6, puf_66_wire_7, puf_66_wire_8,
         puf_67_wire_0, puf_67_wire_1, puf_67_wire_2, puf_67_wire_5, puf_67_wire_6, puf_67_wire_7, puf_67_wire_8, puf_68_wire_0, puf_68_wire_1, puf_68_wire_2, puf_68_wire_5,
         puf_68_wire_6, puf_68_wire_7, puf_68_wire_8, puf_69_wire_0, puf_69_wire_1, puf_69_wire_2, puf_69_wire_5, puf_69_wire_6, puf_69_wire_7, puf_69_wire_8, puf_70_wire_0,
         puf_70_wire_1, puf_70_wire_2, puf_70_wire_5, puf_70_wire_6, puf_70_wire_7, puf_70_wire_8, puf_71_wire_0, puf_71_wire_1, puf_71_wire_2, puf_71_wire_5, puf_71_wire_6,
         puf_71_wire_7, puf_71_wire_8, puf_72_wire_0, puf_72_wire_1, puf_72_wire_2, puf_72_wire_5, puf_72_wire_6, puf_72_wire_7, puf_72_wire_8, puf_73_wire_0, puf_73_wire_1,
         puf_73_wire_2, puf_73_wire_5, puf_73_wire_6, puf_73_wire_7, puf_73_wire_8, puf_74_wire_0, puf_74_wire_1, puf_74_wire_2, puf_74_wire_5, puf_74_wire_6, puf_74_wire_7,
         puf_74_wire_8, puf_75_wire_0, puf_75_wire_1, puf_75_wire_2, puf_75_wire_5, puf_75_wire_6, puf_75_wire_7, puf_75_wire_8, puf_76_wire_0, puf_76_wire_1, puf_76_wire_2,
         puf_76_wire_5, puf_76_wire_6, puf_76_wire_7, puf_76_wire_8, puf_77_wire_0, puf_77_wire_1, puf_77_wire_2, puf_77_wire_5, puf_77_wire_6, puf_77_wire_7, puf_77_wire_8,
         puf_78_wire_0, puf_78_wire_1, puf_78_wire_2, puf_78_wire_5, puf_78_wire_6, puf_78_wire_7, puf_78_wire_8, puf_79_wire_0, puf_79_wire_1, puf_79_wire_2, puf_79_wire_5,
         puf_79_wire_6, puf_79_wire_7, puf_79_wire_8, puf_80_wire_0, puf_80_wire_1, puf_80_wire_2, puf_80_wire_5, puf_80_wire_6, puf_80_wire_7, puf_80_wire_8, puf_81_wire_0,
         puf_81_wire_1, puf_81_wire_2, puf_81_wire_5, puf_81_wire_6, puf_81_wire_7, puf_81_wire_8, puf_82_wire_0, puf_82_wire_1, puf_82_wire_2, puf_82_wire_5, puf_82_wire_6,
         puf_82_wire_7, puf_82_wire_8, puf_83_wire_0, puf_83_wire_1, puf_83_wire_2, puf_83_wire_5, puf_83_wire_6, puf_83_wire_7, puf_83_wire_8, puf_84_wire_0, puf_84_wire_1,
         puf_84_wire_2, puf_84_wire_5, puf_84_wire_6, puf_84_wire_7, puf_84_wire_8, puf_85_wire_0, puf_85_wire_1, puf_85_wire_2, puf_85_wire_5, puf_85_wire_6, puf_85_wire_7,
         puf_85_wire_8, puf_86_wire_0, puf_86_wire_1, puf_86_wire_2, puf_86_wire_5, puf_86_wire_6, puf_86_wire_7, puf_86_wire_8, puf_87_wire_0, puf_87_wire_1, puf_87_wire_2,
         puf_87_wire_5, puf_87_wire_6, puf_87_wire_7, puf_87_wire_8, puf_88_wire_0, puf_88_wire_1, puf_88_wire_2, puf_88_wire_5, puf_88_wire_6, puf_88_wire_7, puf_88_wire_8,
         puf_89_wire_0, puf_89_wire_1, puf_89_wire_2, puf_89_wire_5, puf_89_wire_6, puf_89_wire_7, puf_89_wire_8, puf_90_wire_0, puf_90_wire_1, puf_90_wire_2, puf_90_wire_5,
         puf_90_wire_6, puf_90_wire_7, puf_90_wire_8, puf_91_wire_0, puf_91_wire_1, puf_91_wire_2, puf_91_wire_5, puf_91_wire_6, puf_91_wire_7, puf_91_wire_8, puf_92_wire_0,
         puf_92_wire_1, puf_92_wire_2, puf_92_wire_5, puf_92_wire_6, puf_92_wire_7, puf_92_wire_8, puf_93_wire_0, puf_93_wire_1, puf_93_wire_2, puf_93_wire_5, puf_93_wire_6,
         puf_93_wire_7, puf_93_wire_8, puf_94_wire_0, puf_94_wire_1, puf_94_wire_2, puf_94_wire_5, puf_94_wire_6, puf_94_wire_7, puf_94_wire_8, puf_95_wire_0, puf_95_wire_1,
         puf_95_wire_2, puf_95_wire_5, puf_95_wire_6, puf_95_wire_7, puf_95_wire_8, puf_96_wire_0, puf_96_wire_1, puf_96_wire_2, puf_96_wire_5, puf_96_wire_6, puf_96_wire_7,
         puf_96_wire_8, puf_97_wire_0, puf_97_wire_1, puf_97_wire_2, puf_97_wire_5, puf_97_wire_6, puf_97_wire_7, puf_97_wire_8, puf_98_wire_0, puf_98_wire_1, puf_98_wire_2,
         puf_98_wire_5, puf_98_wire_6, puf_98_wire_7, puf_98_wire_8, puf_99_wire_0, puf_99_wire_1, puf_99_wire_2, puf_99_wire_5, puf_99_wire_6, puf_99_wire_7, puf_99_wire_8,
         puf_100_wire_0, puf_100_wire_1, puf_100_wire_2, puf_100_wire_5, puf_100_wire_6, puf_100_wire_7, puf_100_wire_8, puf_101_wire_0, puf_101_wire_1, puf_101_wire_2, puf_101_wire_5,
         puf_101_wire_6, puf_101_wire_7, puf_101_wire_8, puf_102_wire_0, puf_102_wire_1, puf_102_wire_2, puf_102_wire_5, puf_102_wire_6, puf_102_wire_7, puf_102_wire_8, puf_103_wire_0,
         puf_103_wire_1, puf_103_wire_2, puf_103_wire_5, puf_103_wire_6, puf_103_wire_7, puf_103_wire_8, puf_104_wire_0, puf_104_wire_1, puf_104_wire_2, puf_104_wire_5, puf_104_wire_6,
         puf_104_wire_7, puf_104_wire_8, puf_105_wire_0, puf_105_wire_1, puf_105_wire_2, puf_105_wire_5, puf_105_wire_6, puf_105_wire_7, puf_105_wire_8, puf_106_wire_0, puf_106_wire_1,
         puf_106_wire_2, puf_106_wire_5, puf_106_wire_6, puf_106_wire_7, puf_106_wire_8, puf_107_wire_0, puf_107_wire_1, puf_107_wire_2, puf_107_wire_5, puf_107_wire_6, puf_107_wire_7,
         puf_107_wire_8, puf_108_wire_0, puf_108_wire_1, puf_108_wire_2, puf_108_wire_5, puf_108_wire_6, puf_108_wire_7, puf_108_wire_8, puf_109_wire_0, puf_109_wire_1, puf_109_wire_2,
         puf_109_wire_5, puf_109_wire_6, puf_109_wire_7, puf_109_wire_8, puf_110_wire_0, puf_110_wire_1, puf_110_wire_2, puf_110_wire_5, puf_110_wire_6, puf_110_wire_7, puf_110_wire_8,
         puf_111_wire_0, puf_111_wire_1, puf_111_wire_2, puf_111_wire_5, puf_111_wire_6, puf_111_wire_7, puf_111_wire_8;
    wire [36:5] my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry;
    wire [115:0] my_FIR_filter_firBlock_left_multProducts;
    wire [5:1] inData_in;
    wire [31:0] outData_in;
    wire [31:0] leftOut;
    wire [318:0] my_FIR_filter_firBlock_left_firStep;
    wire [31:0] rightOut;
    wire [31:1] my_FIR_filter_firBlock_right_multProducts;
    wire [33:3] my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry;
    wire [35:7] my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry;
    wire [39:8] my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_220_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_221_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_222_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_223_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_224_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_225_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_226_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_227_carry;
    wire [31:2] my_FIR_filter_firBlock_left_add_228_carry;
    wire [31:2] add_63_carry;


   DFFSR inData_in_reg_31_ ( .CLK(clk),  .D(inData[31]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[36]));
   DFFSR inData_in_reg_30_ ( .CLK(clk),  .D(inData[30]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[115]));
   DFFSR inData_in_reg_29_ ( .CLK(clk),  .D(inData[29]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[114]));
   DFFSR inData_in_reg_28_ ( .CLK(clk),  .D(inData[28]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[113]));
   DFFSR inData_in_reg_27_ ( .CLK(clk),  .D(inData[27]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[112]));
   DFFSR inData_in_reg_26_ ( .CLK(clk),  .D(inData[26]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[111]));
   DFFSR inData_in_reg_25_ ( .CLK(clk),  .D(inData[25]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[110]));
   DFFSR inData_in_reg_24_ ( .CLK(clk),  .D(inData[24]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[109]));
   DFFSR inData_in_reg_23_ ( .CLK(clk),  .D(inData[23]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[108]));
   DFFSR inData_in_reg_22_ ( .CLK(clk),  .D(inData[22]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[107]));
   DFFSR inData_in_reg_21_ ( .CLK(clk),  .D(inData[21]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[106]));
   DFFSR inData_in_reg_20_ ( .CLK(clk),  .D(inData[20]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[105]));
   DFFSR inData_in_reg_19_ ( .CLK(clk),  .D(inData[19]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[104]));
   DFFSR inData_in_reg_18_ ( .CLK(clk),  .D(inData[18]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[103]));
   DFFSR inData_in_reg_17_ ( .CLK(clk),  .D(inData[17]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[102]));
   DFFSR inData_in_reg_16_ ( .CLK(clk),  .D(inData[16]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[101]));
   DFFSR inData_in_reg_15_ ( .CLK(clk),  .D(inData[15]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[100]));
   DFFSR inData_in_reg_14_ ( .CLK(clk),  .D(inData[14]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[99]));
   DFFSR inData_in_reg_13_ ( .CLK(clk),  .D(inData[13]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[98]));
   DFFSR inData_in_reg_12_ ( .CLK(clk),  .D(inData[12]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[97]));
   DFFSR inData_in_reg_11_ ( .CLK(clk),  .D(inData[11]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[96]));
   DFFSR inData_in_reg_10_ ( .CLK(clk),  .D(inData[10]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[95]));
   DFFSR inData_in_reg_9_ ( .CLK(clk),  .D(inData[9]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[94]));
   DFFSR inData_in_reg_8_ ( .CLK(clk),  .D(inData[8]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[93]));
   DFFSR inData_in_reg_7_ ( .CLK(clk),  .D(inData[7]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[92]));
   DFFSR inData_in_reg_6_ ( .CLK(clk),  .D(inData[6]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_multProducts[91]));
   DFFSR inData_in_reg_5_ ( .CLK(clk),  .D(inData[5]),  .R(reset),  .S(VDD), .Q(inData_in[5]));
   DFFSR inData_in_reg_4_ ( .CLK(clk),  .D(inData[4]),  .R(reset),  .S(VDD), .Q(inData_in[4]));
   DFFSR inData_in_reg_3_ ( .CLK(clk),  .D(inData[3]),  .R(reset),  .S(VDD), .Q(inData_in[3]));
   DFFSR inData_in_reg_2_ ( .CLK(clk),  .D(inData[2]),  .R(reset),  .S(VDD), .Q(inData_in[2]));
   DFFSR inData_in_reg_1_ ( .CLK(clk),  .D(inData[1]),  .R(reset),  .S(VDD), .Q(inData_in[1]));
   DFFSR inData_in_reg_0_ ( .CLK(clk),  .D(inData[0]),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_6_));
   DFFSR outData_reg_31_ ( .CLK(clk),  .D(outData_in[31]),  .R(reset),  .S(VDD), .Q(puf_0_wire_1));
   DFFSR outData_reg_30_ ( .CLK(clk),  .D(outData_in[30]),  .R(reset),  .S(VDD), .Q(puf_1_wire_1));
   DFFSR outData_reg_29_ ( .CLK(clk),  .D(outData_in[29]),  .R(reset),  .S(VDD), .Q(puf_2_wire_1));
   DFFSR outData_reg_28_ ( .CLK(clk),  .D(outData_in[28]),  .R(reset),  .S(VDD), .Q(puf_3_wire_1));
   DFFSR outData_reg_27_ ( .CLK(clk),  .D(outData_in[27]),  .R(reset),  .S(VDD), .Q(puf_4_wire_1));
   DFFSR outData_reg_26_ ( .CLK(clk),  .D(outData_in[26]),  .R(reset),  .S(VDD), .Q(puf_5_wire_1));
   DFFSR outData_reg_25_ ( .CLK(clk),  .D(outData_in[25]),  .R(reset),  .S(VDD), .Q(puf_6_wire_1));
   DFFSR outData_reg_24_ ( .CLK(clk),  .D(outData_in[24]),  .R(reset),  .S(VDD), .Q(puf_7_wire_1));
   DFFSR outData_reg_23_ ( .CLK(clk),  .D(outData_in[23]),  .R(reset),  .S(VDD), .Q(puf_8_wire_1));
   DFFSR outData_reg_22_ ( .CLK(clk),  .D(outData_in[22]),  .R(reset),  .S(VDD), .Q(puf_9_wire_1));
   DFFSR outData_reg_21_ ( .CLK(clk),  .D(outData_in[21]),  .R(reset),  .S(VDD), .Q(puf_10_wire_1));
   DFFSR outData_reg_20_ ( .CLK(clk),  .D(outData_in[20]),  .R(reset),  .S(VDD), .Q(puf_11_wire_1));
   DFFSR outData_reg_19_ ( .CLK(clk),  .D(outData_in[19]),  .R(reset),  .S(VDD), .Q(puf_12_wire_1));
   DFFSR outData_reg_18_ ( .CLK(clk),  .D(outData_in[18]),  .R(reset),  .S(VDD), .Q(puf_13_wire_1));
   DFFSR outData_reg_17_ ( .CLK(clk),  .D(outData_in[17]),  .R(reset),  .S(VDD), .Q(puf_14_wire_1));
   DFFSR outData_reg_16_ ( .CLK(clk),  .D(outData_in[16]),  .R(reset),  .S(VDD), .Q(puf_15_wire_1));
   DFFSR outData_reg_15_ ( .CLK(clk),  .D(outData_in[15]),  .R(reset),  .S(VDD), .Q(puf_16_wire_1));
   DFFSR outData_reg_14_ ( .CLK(clk),  .D(outData_in[14]),  .R(reset),  .S(VDD), .Q(puf_17_wire_1));
   DFFSR outData_reg_13_ ( .CLK(clk),  .D(outData_in[13]),  .R(reset),  .S(VDD), .Q(puf_18_wire_1));
   DFFSR outData_reg_12_ ( .CLK(clk),  .D(outData_in[12]),  .R(reset),  .S(VDD), .Q(puf_19_wire_1));
   DFFSR outData_reg_11_ ( .CLK(clk),  .D(outData_in[11]),  .R(reset),  .S(VDD), .Q(puf_20_wire_1));
   DFFSR outData_reg_10_ ( .CLK(clk),  .D(outData_in[10]),  .R(reset),  .S(VDD), .Q(puf_21_wire_1));
   DFFSR outData_reg_9_ ( .CLK(clk),  .D(outData_in[9]),  .R(reset),  .S(VDD), .Q(puf_22_wire_1));
   DFFSR outData_reg_8_ ( .CLK(clk),  .D(outData_in[8]),  .R(reset),  .S(VDD), .Q(puf_23_wire_1));
   DFFSR outData_reg_7_ ( .CLK(clk),  .D(outData_in[7]),  .R(reset),  .S(VDD), .Q(puf_24_wire_1));
   DFFSR outData_reg_6_ ( .CLK(clk),  .D(outData_in[6]),  .R(reset),  .S(VDD), .Q(puf_25_wire_1));
   DFFSR outData_reg_5_ ( .CLK(clk),  .D(outData_in[5]),  .R(reset),  .S(VDD), .Q(puf_26_wire_1));
   DFFSR outData_reg_4_ ( .CLK(clk),  .D(outData_in[4]),  .R(reset),  .S(VDD), .Q(puf_27_wire_1));
   DFFSR outData_reg_3_ ( .CLK(clk),  .D(outData_in[3]),  .R(reset),  .S(VDD), .Q(puf_28_wire_1));
   DFFSR outData_reg_2_ ( .CLK(clk),  .D(outData_in[2]),  .R(reset),  .S(VDD), .Q(puf_29_wire_1));
   DFFSR outData_reg_1_ ( .CLK(clk),  .D(outData_in[1]),  .R(reset),  .S(VDD), .Q(puf_30_wire_1));
   DFFSR outData_reg_0_ ( .CLK(clk),  .D(outData_in[0]),  .R(reset),  .S(VDD), .Q(puf_31_wire_1));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_31_ ( .CLK(clk),  .D(n67),  .R(reset),  .S(VDD), .Q(leftOut[31]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_30_ ( .CLK(clk),  .D(n68),  .R(reset),  .S(VDD), .Q(leftOut[30]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_29_ ( .CLK(clk),  .D(n69),  .R(reset),  .S(VDD), .Q(leftOut[29]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_28_ ( .CLK(clk),  .D(n70),  .R(reset),  .S(VDD), .Q(leftOut[28]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_27_ ( .CLK(clk),  .D(n71),  .R(reset),  .S(VDD), .Q(leftOut[27]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_26_ ( .CLK(clk),  .D(n72),  .R(reset),  .S(VDD), .Q(leftOut[26]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_25_ ( .CLK(clk),  .D(n73),  .R(reset),  .S(VDD), .Q(leftOut[25]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_24_ ( .CLK(clk),  .D(n74),  .R(reset),  .S(VDD), .Q(leftOut[24]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_23_ ( .CLK(clk),  .D(n75),  .R(reset),  .S(VDD), .Q(leftOut[23]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_22_ ( .CLK(clk),  .D(n76),  .R(reset),  .S(VDD), .Q(leftOut[22]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_21_ ( .CLK(clk),  .D(n77),  .R(reset),  .S(VDD), .Q(leftOut[21]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_20_ ( .CLK(clk),  .D(n78),  .R(reset),  .S(VDD), .Q(leftOut[20]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_19_ ( .CLK(clk),  .D(n79),  .R(reset),  .S(VDD), .Q(leftOut[19]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_18_ ( .CLK(clk),  .D(n80),  .R(reset),  .S(VDD), .Q(leftOut[18]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_17_ ( .CLK(clk),  .D(n81),  .R(reset),  .S(VDD), .Q(leftOut[17]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_16_ ( .CLK(clk),  .D(n82),  .R(reset),  .S(VDD), .Q(leftOut[16]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_15_ ( .CLK(clk),  .D(n83),  .R(reset),  .S(VDD), .Q(leftOut[15]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_14_ ( .CLK(clk),  .D(n84),  .R(reset),  .S(VDD), .Q(leftOut[14]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_13_ ( .CLK(clk),  .D(n85),  .R(reset),  .S(VDD), .Q(leftOut[13]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_12_ ( .CLK(clk),  .D(n86),  .R(reset),  .S(VDD), .Q(leftOut[12]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_11_ ( .CLK(clk),  .D(n87),  .R(reset),  .S(VDD), .Q(leftOut[11]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_10_ ( .CLK(clk),  .D(n88),  .R(reset),  .S(VDD), .Q(leftOut[10]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_9_ ( .CLK(clk),  .D(n89),  .R(reset),  .S(VDD), .Q(leftOut[9]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_8_ ( .CLK(clk),  .D(n90),  .R(reset),  .S(VDD), .Q(leftOut[8]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_7_ ( .CLK(clk),  .D(n91),  .R(reset),  .S(VDD), .Q(leftOut[7]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_6_ ( .CLK(clk),  .D(n92),  .R(reset),  .S(VDD), .Q(leftOut[6]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_5_ ( .CLK(clk),  .D(n93),  .R(reset),  .S(VDD), .Q(leftOut[5]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_4_ ( .CLK(clk),  .D(n94),  .R(reset),  .S(VDD), .Q(leftOut[4]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_3_ ( .CLK(clk),  .D(n95),  .R(reset),  .S(VDD), .Q(leftOut[3]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_2_ ( .CLK(clk),  .D(n96),  .R(reset),  .S(VDD), .Q(leftOut[2]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_1_ ( .CLK(clk),  .D(n97),  .R(reset),  .S(VDD), .Q(leftOut[1]));
   DFFSR my_FIR_filter_firBlock_left_Y_reg_0_ ( .CLK(clk),  .D(n98),  .R(reset),  .S(VDD), .Q(leftOut[0]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N257),  .R(reset),  .S(VDD), .Q(puf_32_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N258),  .R(reset),  .S(VDD), .Q(puf_33_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N259),  .R(reset),  .S(VDD), .Q(puf_34_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N260),  .R(reset),  .S(VDD), .Q(puf_35_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N261),  .R(reset),  .S(VDD), .Q(puf_36_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N262),  .R(reset),  .S(VDD), .Q(puf_37_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N263),  .R(reset),  .S(VDD), .Q(puf_38_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N264),  .R(reset),  .S(VDD), .Q(puf_39_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N265),  .R(reset),  .S(VDD), .Q(puf_40_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N266),  .R(reset),  .S(VDD), .Q(puf_41_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N267),  .R(reset),  .S(VDD), .Q(puf_42_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N268),  .R(reset),  .S(VDD), .Q(puf_43_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N269),  .R(reset),  .S(VDD), .Q(puf_44_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N270),  .R(reset),  .S(VDD), .Q(puf_45_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N271),  .R(reset),  .S(VDD), .Q(puf_46_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N272),  .R(reset),  .S(VDD), .Q(puf_47_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N273),  .R(reset),  .S(VDD), .Q(puf_48_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N274),  .R(reset),  .S(VDD), .Q(puf_49_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N275),  .R(reset),  .S(VDD), .Q(puf_50_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N276),  .R(reset),  .S(VDD), .Q(puf_51_wire_1));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N277),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[19]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N278),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[20]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N279),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[21]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N280),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[22]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N281),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[23]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N282),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[24]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N283),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[25]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N284),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[26]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N285),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[27]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N286),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[28]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N287),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[29]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_9__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N288),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[30]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N225),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[31]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N226),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[32]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N227),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[33]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N228),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[34]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N229),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[35]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N230),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[36]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N231),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[37]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N232),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[38]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N233),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[39]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N234),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[40]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N235),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[41]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N236),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[42]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N237),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[43]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N238),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[44]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N239),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[45]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N240),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[46]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N241),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[47]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N242),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[48]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N243),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[49]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N244),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[50]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N245),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[51]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N246),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[52]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N247),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[53]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N248),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[54]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N249),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[55]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N250),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[56]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N251),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[57]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N252),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[58]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N253),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[59]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N254),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[60]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N255),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[61]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_8__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N256),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[62]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N193),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[63]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N194),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[64]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N195),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[65]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N196),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[66]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N197),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[67]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N198),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[68]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N199),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[69]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N200),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[70]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N201),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[71]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N202),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[72]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N203),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[73]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N204),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[74]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N205),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[75]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N206),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[76]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N207),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[77]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N208),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[78]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N209),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[79]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N210),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[80]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N211),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[81]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N212),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[82]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N213),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[83]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N214),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[84]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N215),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[85]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N216),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[86]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N217),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[87]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N218),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[88]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N219),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[89]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N220),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[90]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N221),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[91]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N222),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[92]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N223),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[93]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_7__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N224),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[94]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N161),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[95]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N162),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[96]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N163),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[97]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N164),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[98]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N165),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[99]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N166),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[100]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N167),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[101]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N168),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[102]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N169),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[103]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N170),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[104]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N171),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[105]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N172),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[106]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N173),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[107]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N174),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[108]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N175),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[109]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N176),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[110]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N177),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[111]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N178),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[112]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N179),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[113]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N180),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[114]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N181),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[115]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N182),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[116]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N183),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[117]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N184),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[118]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N185),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[119]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N186),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[120]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N187),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[121]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N188),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[122]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N189),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[123]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N190),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[124]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N191),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[125]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_6__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N192),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[126]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N129),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[127]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N130),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[128]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N131),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[129]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N132),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[130]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N133),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[131]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N134),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[132]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N135),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[133]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N136),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[134]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N137),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[135]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N138),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[136]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N139),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[137]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N140),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[138]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N141),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[139]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N142),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[140]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N143),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[141]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N144),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[142]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N145),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[143]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N146),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[144]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N147),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[145]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N148),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[146]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N149),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[147]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N150),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[148]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N151),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[149]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N152),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[150]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N153),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[151]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N154),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[152]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N155),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[153]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N156),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[154]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N157),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[155]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N158),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[156]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N159),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[157]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_5__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N160),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[158]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N97),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[159]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N98),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[160]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N99),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[161]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N100),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[162]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N101),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[163]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N102),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[164]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N103),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[165]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N104),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[166]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N105),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[167]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N106),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[168]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N107),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[169]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N108),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[170]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N109),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[171]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N110),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[172]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N111),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[173]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N112),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[174]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N113),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[175]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N114),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[176]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N115),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[177]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N116),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[178]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N117),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[179]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N118),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[180]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N119),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[181]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N120),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[182]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N121),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[183]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N122),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[184]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N123),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[185]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N124),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[186]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N125),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[187]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N126),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[188]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N127),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[189]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_4__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N128),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[190]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N65),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[191]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N66),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[192]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N67),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[193]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N68),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[194]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N69),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[195]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N70),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[196]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N71),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[197]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N72),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[198]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N73),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[199]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N74),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[200]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N75),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[201]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N76),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[202]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N77),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[203]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N78),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[204]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N79),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[205]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N80),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[206]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N81),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[207]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N82),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[208]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N83),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[209]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N84),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[210]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N85),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[211]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N86),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[212]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N87),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[213]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N88),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[214]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N89),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[215]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N90),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[216]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N91),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[217]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N92),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[218]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N93),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[219]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N94),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[220]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N95),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[221]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_3__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N96),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[222]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N33),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[223]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N34),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[224]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N35),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[225]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N36),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[226]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N37),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[227]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N38),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[228]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N39),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[229]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N40),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[230]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N41),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[231]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N42),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[232]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N43),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[233]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N44),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[234]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N45),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[235]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N46),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[236]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N47),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[237]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N48),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[238]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N49),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[239]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N50),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[240]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N51),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[241]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N52),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[242]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N53),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[243]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N54),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[244]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N55),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[245]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N56),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[246]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N57),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[247]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N58),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[248]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N59),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[249]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N60),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[250]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N61),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[251]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N62),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[252]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N63),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[253]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_2__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N64),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[254]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__0_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N1),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[255]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N2),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[256]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N3),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[257]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N4),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[258]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N5),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[259]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N6),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[260]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N7),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[261]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N8),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[262]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N9),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[263]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N10),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[264]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N11),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[265]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N12),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[266]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N13),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[267]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N14),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[268]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N15),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[269]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N16),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[270]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N17),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[271]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N18),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[272]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N19),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[273]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N20),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[274]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N21),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[275]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N22),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[276]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N23),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[277]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N24),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[278]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N25),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[279]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N26),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[280]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N27),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[281]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N28),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[282]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N29),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[283]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N30),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[284]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N31),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[285]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_1__31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_left_N32),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[286]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__0_ ( .CLK(clk),  .D(n317),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[287]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__1_ ( .CLK(clk),  .D(n485),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[288]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__2_ ( .CLK(clk),  .D(n483),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[289]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__3_ ( .CLK(clk),  .D(n484),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[290]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__4_ ( .CLK(clk),  .D(n482),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[291]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__5_ ( .CLK(clk),  .D(n316),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[292]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__6_ ( .CLK(clk),  .D(n315),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[293]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__7_ ( .CLK(clk),  .D(n314),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[294]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__8_ ( .CLK(clk),  .D(n313),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[295]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__9_ ( .CLK(clk),  .D(n481),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[296]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__10_ ( .CLK(clk),  .D(n480),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[297]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__11_ ( .CLK(clk),  .D(n479),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[298]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__12_ ( .CLK(clk),  .D(n478),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[299]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__13_ ( .CLK(clk),  .D(n312),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[300]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__14_ ( .CLK(clk),  .D(n311),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[301]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__15_ ( .CLK(clk),  .D(n310),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[302]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__16_ ( .CLK(clk),  .D(n309),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[303]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__17_ ( .CLK(clk),  .D(n477),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[304]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__18_ ( .CLK(clk),  .D(n476),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[305]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__19_ ( .CLK(clk),  .D(n475),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[306]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__20_ ( .CLK(clk),  .D(n474),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[307]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__21_ ( .CLK(clk),  .D(n308),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[308]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__22_ ( .CLK(clk),  .D(n307),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[309]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__23_ ( .CLK(clk),  .D(n306),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[310]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__24_ ( .CLK(clk),  .D(n305),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[311]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__25_ ( .CLK(clk),  .D(n486),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[312]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__26_ ( .CLK(clk),  .D(n486),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[313]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__27_ ( .CLK(clk),  .D(n486),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[314]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__28_ ( .CLK(clk),  .D(n486),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[315]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__29_ ( .CLK(clk),  .D(n486),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[316]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__30_ ( .CLK(clk),  .D(n486),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[317]));
   DFFSR my_FIR_filter_firBlock_left_firStep_reg_0__31_ ( .CLK(clk),  .D(n486),  .R(reset),  .S(VDD), .Q(my_FIR_filter_firBlock_left_firStep[318]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_0_ ( .CLK(clk),  .D(outData_in[0]),  .R(reset),  .S(VDD), .Q(rightOut[0]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_1_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[1]),  .R(reset),  .S(VDD), .Q(rightOut[1]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_2_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[2]),  .R(reset),  .S(VDD), .Q(rightOut[2]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_3_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[3]),  .R(reset),  .S(VDD), .Q(rightOut[3]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_4_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[4]),  .R(reset),  .S(VDD), .Q(rightOut[4]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_5_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[5]),  .R(reset),  .S(VDD), .Q(rightOut[5]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_6_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[6]),  .R(reset),  .S(VDD), .Q(rightOut[6]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_7_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[7]),  .R(reset),  .S(VDD), .Q(rightOut[7]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_8_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[8]),  .R(reset),  .S(VDD), .Q(rightOut[8]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_9_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[9]),  .R(reset),  .S(VDD), .Q(rightOut[9]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_10_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[10]),  .R(reset),  .S(VDD), .Q(rightOut[10]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_11_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[11]),  .R(reset),  .S(VDD), .Q(rightOut[11]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_12_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[12]),  .R(reset),  .S(VDD), .Q(rightOut[12]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_13_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[13]),  .R(reset),  .S(VDD), .Q(rightOut[13]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_14_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[14]),  .R(reset),  .S(VDD), .Q(rightOut[14]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_15_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[15]),  .R(reset),  .S(VDD), .Q(rightOut[15]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_16_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[16]),  .R(reset),  .S(VDD), .Q(rightOut[16]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_17_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[17]),  .R(reset),  .S(VDD), .Q(rightOut[17]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_18_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[18]),  .R(reset),  .S(VDD), .Q(rightOut[18]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_19_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[19]),  .R(reset),  .S(VDD), .Q(rightOut[19]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_20_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[20]),  .R(reset),  .S(VDD), .Q(rightOut[20]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_21_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[21]),  .R(reset),  .S(VDD), .Q(rightOut[21]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_22_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[22]),  .R(reset),  .S(VDD), .Q(rightOut[22]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_23_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[23]),  .R(reset),  .S(VDD), .Q(rightOut[23]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_24_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[24]),  .R(reset),  .S(VDD), .Q(rightOut[24]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_25_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[25]),  .R(reset),  .S(VDD), .Q(rightOut[25]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_26_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[26]),  .R(reset),  .S(VDD), .Q(rightOut[26]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_27_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[27]),  .R(reset),  .S(VDD), .Q(rightOut[27]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_28_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[28]),  .R(reset),  .S(VDD), .Q(rightOut[28]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_29_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[29]),  .R(reset),  .S(VDD), .Q(rightOut[29]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_30_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[30]),  .R(reset),  .S(VDD), .Q(rightOut[30]));
   DFFSR my_FIR_filter_firBlock_right_Y_reg_31_ ( .CLK(clk),  .D(my_FIR_filter_firBlock_right_multProducts[31]),  .R(reset),  .S(VDD), .Q(rightOut[31]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_2 ( .A(n103),  .B(n571),  .C(n517), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[3]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_8_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_3 ( .A(n137),  .B(n570),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[3]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[4]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_9_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_4 ( .A(n473),  .B(n569),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[4]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[5]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_10_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_5 ( .A(n303),  .B(n568),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[5]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[6]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_11_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_6 ( .A(n138),  .B(n567),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[6]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[7]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_12_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_7 ( .A(n304),  .B(n566),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[7]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[8]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_13_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_8 ( .A(n317),  .B(n565),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[8]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[9]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_14_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_9 ( .A(n485),  .B(n564),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[9]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[10]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_15_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_10 ( .A(n483),  .B(n563),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[10]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[11]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_16_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_11 ( .A(n484),  .B(n562),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[11]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[12]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_17_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_12 ( .A(n482),  .B(n561),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[12]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[13]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_18_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_13 ( .A(n316),  .B(n560),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[13]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[14]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_19_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_14 ( .A(n315),  .B(n559),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[14]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[15]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_20_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_15 ( .A(n314),  .B(n558),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[15]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[16]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_21_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_16 ( .A(n313),  .B(n557),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[16]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[17]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_22_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_17 ( .A(n481),  .B(n556),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[17]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[18]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_23_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_18 ( .A(n480),  .B(n555),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[18]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[19]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_24_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_19 ( .A(n479),  .B(n554),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[19]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[20]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_25_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_20 ( .A(n478),  .B(n553),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[20]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[21]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_26_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_21 ( .A(n312),  .B(n552),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[21]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[22]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_27_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_22 ( .A(n311),  .B(n551),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[22]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[23]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_28_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_23 ( .A(n310),  .B(n550),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[23]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[24]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_29_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_24 ( .A(n309),  .B(n549),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[24]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[25]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_30_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_25 ( .A(n477),  .B(n548),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[25]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[26]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_31_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_26 ( .A(n476),  .B(n547),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[26]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[27]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_32_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_27 ( .A(n475),  .B(n546),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[27]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[28]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_33_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_28 ( .A(n474),  .B(n545),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[28]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[29]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_34_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_29 ( .A(n308),  .B(n544),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[29]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[30]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_35_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_30 ( .A(n307),  .B(n543),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[30]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[31]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_36_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_31 ( .A(n306),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[31]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[32]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_37_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_U2_32 ( .A(n305),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[32]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[33]), .YS(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_38_));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_7 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_13_),  .B(n138),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[7]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[8]), .YS(my_FIR_filter_firBlock_left_multProducts[62]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_8 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_14_),  .B(n304),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[8]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[9]), .YS(my_FIR_filter_firBlock_left_multProducts[63]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_9 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_15_),  .B(n317),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[9]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[10]), .YS(my_FIR_filter_firBlock_left_multProducts[64]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_10 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_16_),  .B(n485),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[10]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[11]), .YS(my_FIR_filter_firBlock_left_multProducts[65]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_11 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_17_),  .B(n483),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[11]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[12]), .YS(my_FIR_filter_firBlock_left_multProducts[66]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_12 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_18_),  .B(n484),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[12]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[13]), .YS(my_FIR_filter_firBlock_left_multProducts[67]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_13 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_19_),  .B(n482),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[13]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[14]), .YS(my_FIR_filter_firBlock_left_multProducts[68]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_14 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_20_),  .B(n316),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[14]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[15]), .YS(my_FIR_filter_firBlock_left_multProducts[69]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_15 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_21_),  .B(n315),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[15]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[16]), .YS(my_FIR_filter_firBlock_left_multProducts[70]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_16 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_22_),  .B(n314),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[16]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[17]), .YS(my_FIR_filter_firBlock_left_multProducts[71]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_17 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_23_),  .B(n313),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[17]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[18]), .YS(my_FIR_filter_firBlock_left_multProducts[72]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_18 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_24_),  .B(n481),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[18]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[19]), .YS(my_FIR_filter_firBlock_left_multProducts[73]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_19 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_25_),  .B(n480),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[19]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[20]), .YS(my_FIR_filter_firBlock_left_multProducts[74]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_20 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_26_),  .B(n479),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[20]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[21]), .YS(my_FIR_filter_firBlock_left_multProducts[75]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_21 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_27_),  .B(n478),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[21]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[22]), .YS(my_FIR_filter_firBlock_left_multProducts[76]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_22 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_28_),  .B(n312),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[22]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[23]), .YS(my_FIR_filter_firBlock_left_multProducts[77]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_23 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_29_),  .B(n311),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[23]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[24]), .YS(my_FIR_filter_firBlock_left_multProducts[78]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_24 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_30_),  .B(n310),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[24]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[25]), .YS(my_FIR_filter_firBlock_left_multProducts[79]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_25 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_31_),  .B(n309),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[25]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[26]), .YS(my_FIR_filter_firBlock_left_multProducts[80]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_26 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_32_),  .B(n477),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[26]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[27]), .YS(my_FIR_filter_firBlock_left_multProducts[81]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_27 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_33_),  .B(n476),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[27]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[28]), .YS(my_FIR_filter_firBlock_left_multProducts[82]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_28 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_34_),  .B(n475),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[28]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[29]), .YS(my_FIR_filter_firBlock_left_multProducts[83]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_29 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_35_),  .B(n474),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[29]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[30]), .YS(my_FIR_filter_firBlock_left_multProducts[84]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_30 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_36_),  .B(n308),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[30]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[31]), .YS(my_FIR_filter_firBlock_left_multProducts[85]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_31 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_37_),  .B(n307),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[31]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[32]), .YS(my_FIR_filter_firBlock_left_multProducts[86]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_32 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_38_),  .B(n306),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[32]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[33]), .YS(my_FIR_filter_firBlock_left_multProducts[87]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_33 ( .A(n541),  .B(n305),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[33]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[34]), .YS(my_FIR_filter_firBlock_left_multProducts[88]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_34 ( .A(n541),  .B(n486),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[34]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[35]), .YS(my_FIR_filter_firBlock_left_multProducts[89]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_U1_35 ( .A(n541),  .B(n486),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[35]), .YS(my_FIR_filter_firBlock_left_multProducts[90]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_5 ( .A(n304),  .B(n137),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[5]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[6]), .YS(my_FIR_filter_firBlock_left_multProducts[32]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_6 ( .A(n317),  .B(n473),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[6]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[7]), .YS(my_FIR_filter_firBlock_left_multProducts[33]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_7 ( .A(n485),  .B(n303),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[7]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[8]), .YS(my_FIR_filter_firBlock_left_multProducts[34]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_8 ( .A(n483),  .B(n138),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[8]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[9]), .YS(my_FIR_filter_firBlock_left_multProducts[35]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_9 ( .A(n484),  .B(n304),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[9]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[10]), .YS(my_FIR_filter_firBlock_left_multProducts[36]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_10 ( .A(n482),  .B(n317),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[10]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[11]), .YS(my_FIR_filter_firBlock_left_multProducts[37]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_11 ( .A(n316),  .B(n485),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[11]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[12]), .YS(my_FIR_filter_firBlock_left_multProducts[38]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_12 ( .A(n315),  .B(n483),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[12]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[13]), .YS(my_FIR_filter_firBlock_left_multProducts[39]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_13 ( .A(n314),  .B(n484),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[13]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[14]), .YS(my_FIR_filter_firBlock_left_multProducts[40]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_14 ( .A(n313),  .B(n482),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[14]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[15]), .YS(my_FIR_filter_firBlock_left_multProducts[41]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_15 ( .A(n481),  .B(n316),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[15]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[16]), .YS(my_FIR_filter_firBlock_left_multProducts[42]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_16 ( .A(n480),  .B(n315),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[16]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[17]), .YS(my_FIR_filter_firBlock_left_multProducts[43]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_17 ( .A(n479),  .B(n314),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[17]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[18]), .YS(my_FIR_filter_firBlock_left_multProducts[44]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_18 ( .A(n478),  .B(n313),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[18]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[19]), .YS(my_FIR_filter_firBlock_left_multProducts[45]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_19 ( .A(n312),  .B(n481),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[19]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[20]), .YS(my_FIR_filter_firBlock_left_multProducts[46]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_20 ( .A(n311),  .B(n480),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[20]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[21]), .YS(my_FIR_filter_firBlock_left_multProducts[47]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_21 ( .A(n310),  .B(n479),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[21]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[22]), .YS(my_FIR_filter_firBlock_left_multProducts[48]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_22 ( .A(n309),  .B(n478),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[22]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[23]), .YS(my_FIR_filter_firBlock_left_multProducts[49]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_23 ( .A(n477),  .B(n312),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[23]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[24]), .YS(my_FIR_filter_firBlock_left_multProducts[50]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_24 ( .A(n476),  .B(n311),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[24]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[25]), .YS(my_FIR_filter_firBlock_left_multProducts[51]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_25 ( .A(n475),  .B(n310),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[25]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[26]), .YS(my_FIR_filter_firBlock_left_multProducts[52]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_26 ( .A(n474),  .B(n309),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[26]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[27]), .YS(my_FIR_filter_firBlock_left_multProducts[53]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_27 ( .A(n308),  .B(n477),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[27]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[28]), .YS(my_FIR_filter_firBlock_left_multProducts[54]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_28 ( .A(n307),  .B(n476),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[28]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[29]), .YS(my_FIR_filter_firBlock_left_multProducts[55]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_29 ( .A(n306),  .B(n475),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[29]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[30]), .YS(my_FIR_filter_firBlock_left_multProducts[56]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_30 ( .A(n305),  .B(n474),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[30]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[31]), .YS(my_FIR_filter_firBlock_left_multProducts[57]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_31 ( .A(n486),  .B(n308),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[31]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[32]), .YS(my_FIR_filter_firBlock_left_multProducts[58]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_32 ( .A(n486),  .B(n307),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[32]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[33]), .YS(my_FIR_filter_firBlock_left_multProducts[59]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_33 ( .A(n486),  .B(n306),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[33]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[34]), .YS(my_FIR_filter_firBlock_left_multProducts[60]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_U1_34 ( .A(n486),  .B(n305),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[34]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[35]), .YS(my_FIR_filter_firBlock_left_multProducts[61]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_8 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_8_),  .B(n565),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[8]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[9]), .YS(my_FIR_filter_firBlock_left_multProducts[0]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_9 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_9_),  .B(n564),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[9]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[10]), .YS(my_FIR_filter_firBlock_left_multProducts[1]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_10 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_10_),  .B(n563),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[10]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[11]), .YS(my_FIR_filter_firBlock_left_multProducts[2]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_11 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_11_),  .B(n562),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[11]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[12]), .YS(my_FIR_filter_firBlock_left_multProducts[3]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_12 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_12_),  .B(n561),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[12]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[13]), .YS(my_FIR_filter_firBlock_left_multProducts[4]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_13 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_13_),  .B(n560),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[13]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[14]), .YS(my_FIR_filter_firBlock_left_multProducts[5]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_14 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_14_),  .B(n559),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[14]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[15]), .YS(my_FIR_filter_firBlock_left_multProducts[6]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_15 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_15_),  .B(n558),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[15]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[16]), .YS(my_FIR_filter_firBlock_left_multProducts[7]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_16 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_16_),  .B(n557),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[16]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[17]), .YS(my_FIR_filter_firBlock_left_multProducts[8]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_17 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_17_),  .B(n556),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[17]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[18]), .YS(my_FIR_filter_firBlock_left_multProducts[9]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_18 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_18_),  .B(n555),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[18]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[19]), .YS(my_FIR_filter_firBlock_left_multProducts[10]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_19 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_19_),  .B(n554),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[19]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[20]), .YS(my_FIR_filter_firBlock_left_multProducts[11]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_20 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_20_),  .B(n553),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[20]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[21]), .YS(my_FIR_filter_firBlock_left_multProducts[12]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_21 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_21_),  .B(n552),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[21]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[22]), .YS(my_FIR_filter_firBlock_left_multProducts[13]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_22 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_22_),  .B(n551),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[22]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[23]), .YS(my_FIR_filter_firBlock_left_multProducts[14]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_23 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_23_),  .B(n550),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[23]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[24]), .YS(my_FIR_filter_firBlock_left_multProducts[15]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_24 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_24_),  .B(n549),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[24]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[25]), .YS(my_FIR_filter_firBlock_left_multProducts[16]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_25 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_25_),  .B(n548),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[25]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[26]), .YS(my_FIR_filter_firBlock_left_multProducts[17]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_26 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_26_),  .B(n547),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[26]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[27]), .YS(my_FIR_filter_firBlock_left_multProducts[18]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_27 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_27_),  .B(n546),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[27]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[28]), .YS(my_FIR_filter_firBlock_left_multProducts[19]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_28 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_28_),  .B(n545),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[28]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[29]), .YS(my_FIR_filter_firBlock_left_multProducts[20]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_29 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_29_),  .B(n544),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[29]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[30]), .YS(my_FIR_filter_firBlock_left_multProducts[21]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_30 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_30_),  .B(n543),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[30]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[31]), .YS(my_FIR_filter_firBlock_left_multProducts[22]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_31 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_31_),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[31]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[32]), .YS(my_FIR_filter_firBlock_left_multProducts[23]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_32 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_32_),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[32]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[33]), .YS(my_FIR_filter_firBlock_left_multProducts[24]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_33 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_33_),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[33]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[34]), .YS(my_FIR_filter_firBlock_left_multProducts[25]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_34 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_34_),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[34]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[35]), .YS(my_FIR_filter_firBlock_left_multProducts[26]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_35 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_35_),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[35]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[36]), .YS(my_FIR_filter_firBlock_left_multProducts[27]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_36 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_36_),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[36]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[37]), .YS(my_FIR_filter_firBlock_left_multProducts[28]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_37 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_37_),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[37]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[38]), .YS(my_FIR_filter_firBlock_left_multProducts[29]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_38 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_38_),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[38]), .YC(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[39]), .YS(my_FIR_filter_firBlock_left_multProducts[30]));
   FAX1 my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_U2_39 ( .A(n541),  .B(n542),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[39]), .YS(my_FIR_filter_firBlock_left_multProducts[31]));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_1 ( .A(n298),  .B(my_FIR_filter_firBlock_left_multProducts[63]),  .C(n518), .YC(my_FIR_filter_firBlock_left_add_220_carry[2]), .YS(my_FIR_filter_firBlock_left_N2));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_2 ( .A(n276),  .B(my_FIR_filter_firBlock_left_multProducts[64]),  .C(my_FIR_filter_firBlock_left_add_220_carry[2]), .YC(my_FIR_filter_firBlock_left_add_220_carry[3]), .YS(my_FIR_filter_firBlock_left_N3));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_3 ( .A(n277),  .B(my_FIR_filter_firBlock_left_multProducts[65]),  .C(my_FIR_filter_firBlock_left_add_220_carry[3]), .YC(my_FIR_filter_firBlock_left_add_220_carry[4]), .YS(my_FIR_filter_firBlock_left_N4));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_4 ( .A(n278),  .B(my_FIR_filter_firBlock_left_multProducts[66]),  .C(my_FIR_filter_firBlock_left_add_220_carry[4]), .YC(my_FIR_filter_firBlock_left_add_220_carry[5]), .YS(my_FIR_filter_firBlock_left_N5));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_5 ( .A(n123),  .B(my_FIR_filter_firBlock_left_multProducts[67]),  .C(my_FIR_filter_firBlock_left_add_220_carry[5]), .YC(my_FIR_filter_firBlock_left_add_220_carry[6]), .YS(my_FIR_filter_firBlock_left_N6));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_6 ( .A(n124),  .B(my_FIR_filter_firBlock_left_multProducts[68]),  .C(my_FIR_filter_firBlock_left_add_220_carry[6]), .YC(my_FIR_filter_firBlock_left_add_220_carry[7]), .YS(my_FIR_filter_firBlock_left_N7));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_7 ( .A(n125),  .B(my_FIR_filter_firBlock_left_multProducts[69]),  .C(my_FIR_filter_firBlock_left_add_220_carry[7]), .YC(my_FIR_filter_firBlock_left_add_220_carry[8]), .YS(my_FIR_filter_firBlock_left_N8));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_8 ( .A(n126),  .B(my_FIR_filter_firBlock_left_multProducts[70]),  .C(my_FIR_filter_firBlock_left_add_220_carry[8]), .YC(my_FIR_filter_firBlock_left_add_220_carry[9]), .YS(my_FIR_filter_firBlock_left_N9));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_9 ( .A(n279),  .B(my_FIR_filter_firBlock_left_multProducts[71]),  .C(my_FIR_filter_firBlock_left_add_220_carry[9]), .YC(my_FIR_filter_firBlock_left_add_220_carry[10]), .YS(my_FIR_filter_firBlock_left_N10));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_10 ( .A(n280),  .B(my_FIR_filter_firBlock_left_multProducts[72]),  .C(my_FIR_filter_firBlock_left_add_220_carry[10]), .YC(my_FIR_filter_firBlock_left_add_220_carry[11]), .YS(my_FIR_filter_firBlock_left_N11));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_11 ( .A(n281),  .B(my_FIR_filter_firBlock_left_multProducts[73]),  .C(my_FIR_filter_firBlock_left_add_220_carry[11]), .YC(my_FIR_filter_firBlock_left_add_220_carry[12]), .YS(my_FIR_filter_firBlock_left_N12));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_12 ( .A(n282),  .B(my_FIR_filter_firBlock_left_multProducts[74]),  .C(my_FIR_filter_firBlock_left_add_220_carry[12]), .YC(my_FIR_filter_firBlock_left_add_220_carry[13]), .YS(my_FIR_filter_firBlock_left_N13));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_13 ( .A(n127),  .B(my_FIR_filter_firBlock_left_multProducts[75]),  .C(my_FIR_filter_firBlock_left_add_220_carry[13]), .YC(my_FIR_filter_firBlock_left_add_220_carry[14]), .YS(my_FIR_filter_firBlock_left_N14));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_14 ( .A(n128),  .B(my_FIR_filter_firBlock_left_multProducts[76]),  .C(my_FIR_filter_firBlock_left_add_220_carry[14]), .YC(my_FIR_filter_firBlock_left_add_220_carry[15]), .YS(my_FIR_filter_firBlock_left_N15));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_15 ( .A(n129),  .B(my_FIR_filter_firBlock_left_multProducts[77]),  .C(my_FIR_filter_firBlock_left_add_220_carry[15]), .YC(my_FIR_filter_firBlock_left_add_220_carry[16]), .YS(my_FIR_filter_firBlock_left_N16));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_16 ( .A(n130),  .B(my_FIR_filter_firBlock_left_multProducts[78]),  .C(my_FIR_filter_firBlock_left_add_220_carry[16]), .YC(my_FIR_filter_firBlock_left_add_220_carry[17]), .YS(my_FIR_filter_firBlock_left_N17));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_17 ( .A(n283),  .B(my_FIR_filter_firBlock_left_multProducts[79]),  .C(my_FIR_filter_firBlock_left_add_220_carry[17]), .YC(my_FIR_filter_firBlock_left_add_220_carry[18]), .YS(my_FIR_filter_firBlock_left_N18));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_18 ( .A(n284),  .B(my_FIR_filter_firBlock_left_multProducts[80]),  .C(my_FIR_filter_firBlock_left_add_220_carry[18]), .YC(my_FIR_filter_firBlock_left_add_220_carry[19]), .YS(my_FIR_filter_firBlock_left_N19));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_19 ( .A(n285),  .B(my_FIR_filter_firBlock_left_multProducts[81]),  .C(my_FIR_filter_firBlock_left_add_220_carry[19]), .YC(my_FIR_filter_firBlock_left_add_220_carry[20]), .YS(my_FIR_filter_firBlock_left_N20));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_20 ( .A(n286),  .B(my_FIR_filter_firBlock_left_multProducts[82]),  .C(my_FIR_filter_firBlock_left_add_220_carry[20]), .YC(my_FIR_filter_firBlock_left_add_220_carry[21]), .YS(my_FIR_filter_firBlock_left_N21));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_21 ( .A(n131),  .B(my_FIR_filter_firBlock_left_multProducts[83]),  .C(my_FIR_filter_firBlock_left_add_220_carry[21]), .YC(my_FIR_filter_firBlock_left_add_220_carry[22]), .YS(my_FIR_filter_firBlock_left_N22));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_22 ( .A(n132),  .B(my_FIR_filter_firBlock_left_multProducts[84]),  .C(my_FIR_filter_firBlock_left_add_220_carry[22]), .YC(my_FIR_filter_firBlock_left_add_220_carry[23]), .YS(my_FIR_filter_firBlock_left_N23));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_23 ( .A(n133),  .B(my_FIR_filter_firBlock_left_multProducts[85]),  .C(my_FIR_filter_firBlock_left_add_220_carry[23]), .YC(my_FIR_filter_firBlock_left_add_220_carry[24]), .YS(my_FIR_filter_firBlock_left_N24));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_24 ( .A(n134),  .B(my_FIR_filter_firBlock_left_multProducts[86]),  .C(my_FIR_filter_firBlock_left_add_220_carry[24]), .YC(my_FIR_filter_firBlock_left_add_220_carry[25]), .YS(my_FIR_filter_firBlock_left_N25));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_25 ( .A(n287),  .B(my_FIR_filter_firBlock_left_multProducts[87]),  .C(my_FIR_filter_firBlock_left_add_220_carry[25]), .YC(my_FIR_filter_firBlock_left_add_220_carry[26]), .YS(my_FIR_filter_firBlock_left_N26));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_26 ( .A(n288),  .B(my_FIR_filter_firBlock_left_multProducts[88]),  .C(my_FIR_filter_firBlock_left_add_220_carry[26]), .YC(my_FIR_filter_firBlock_left_add_220_carry[27]), .YS(my_FIR_filter_firBlock_left_N27));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_27 ( .A(n289),  .B(my_FIR_filter_firBlock_left_multProducts[89]),  .C(my_FIR_filter_firBlock_left_add_220_carry[27]), .YC(my_FIR_filter_firBlock_left_add_220_carry[28]), .YS(my_FIR_filter_firBlock_left_N28));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_28 ( .A(n290),  .B(my_FIR_filter_firBlock_left_multProducts[90]),  .C(my_FIR_filter_firBlock_left_add_220_carry[28]), .YC(my_FIR_filter_firBlock_left_add_220_carry[29]), .YS(my_FIR_filter_firBlock_left_N29));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_29 ( .A(n291),  .B(my_FIR_filter_firBlock_left_multProducts[90]),  .C(my_FIR_filter_firBlock_left_add_220_carry[29]), .YC(my_FIR_filter_firBlock_left_add_220_carry[30]), .YS(my_FIR_filter_firBlock_left_N30));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_30 ( .A(n292),  .B(my_FIR_filter_firBlock_left_multProducts[90]),  .C(my_FIR_filter_firBlock_left_add_220_carry[30]), .YC(my_FIR_filter_firBlock_left_add_220_carry[31]), .YS(my_FIR_filter_firBlock_left_N31));
   FAX1 my_FIR_filter_firBlock_left_add_220_U1_31 ( .A(n293),  .B(my_FIR_filter_firBlock_left_multProducts[90]),  .C(my_FIR_filter_firBlock_left_add_220_carry[31]), .YS(my_FIR_filter_firBlock_left_N32));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_1 ( .A(n467),  .B(my_FIR_filter_firBlock_left_multProducts[34]),  .C(n519), .YC(my_FIR_filter_firBlock_left_add_221_carry[2]), .YS(my_FIR_filter_firBlock_left_N34));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_2 ( .A(n432),  .B(my_FIR_filter_firBlock_left_multProducts[35]),  .C(my_FIR_filter_firBlock_left_add_221_carry[2]), .YC(my_FIR_filter_firBlock_left_add_221_carry[3]), .YS(my_FIR_filter_firBlock_left_N35));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_3 ( .A(n433),  .B(my_FIR_filter_firBlock_left_multProducts[36]),  .C(my_FIR_filter_firBlock_left_add_221_carry[3]), .YC(my_FIR_filter_firBlock_left_add_221_carry[4]), .YS(my_FIR_filter_firBlock_left_N36));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_4 ( .A(n434),  .B(my_FIR_filter_firBlock_left_multProducts[37]),  .C(my_FIR_filter_firBlock_left_add_221_carry[4]), .YC(my_FIR_filter_firBlock_left_add_221_carry[5]), .YS(my_FIR_filter_firBlock_left_N37));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_5 ( .A(n435),  .B(my_FIR_filter_firBlock_left_multProducts[38]),  .C(my_FIR_filter_firBlock_left_add_221_carry[5]), .YC(my_FIR_filter_firBlock_left_add_221_carry[6]), .YS(my_FIR_filter_firBlock_left_N38));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_6 ( .A(n436),  .B(my_FIR_filter_firBlock_left_multProducts[39]),  .C(my_FIR_filter_firBlock_left_add_221_carry[6]), .YC(my_FIR_filter_firBlock_left_add_221_carry[7]), .YS(my_FIR_filter_firBlock_left_N39));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_7 ( .A(n437),  .B(my_FIR_filter_firBlock_left_multProducts[40]),  .C(my_FIR_filter_firBlock_left_add_221_carry[7]), .YC(my_FIR_filter_firBlock_left_add_221_carry[8]), .YS(my_FIR_filter_firBlock_left_N40));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_8 ( .A(n438),  .B(my_FIR_filter_firBlock_left_multProducts[41]),  .C(my_FIR_filter_firBlock_left_add_221_carry[8]), .YC(my_FIR_filter_firBlock_left_add_221_carry[9]), .YS(my_FIR_filter_firBlock_left_N41));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_9 ( .A(n439),  .B(my_FIR_filter_firBlock_left_multProducts[42]),  .C(my_FIR_filter_firBlock_left_add_221_carry[9]), .YC(my_FIR_filter_firBlock_left_add_221_carry[10]), .YS(my_FIR_filter_firBlock_left_N42));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_10 ( .A(n440),  .B(my_FIR_filter_firBlock_left_multProducts[43]),  .C(my_FIR_filter_firBlock_left_add_221_carry[10]), .YC(my_FIR_filter_firBlock_left_add_221_carry[11]), .YS(my_FIR_filter_firBlock_left_N43));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_11 ( .A(n441),  .B(my_FIR_filter_firBlock_left_multProducts[44]),  .C(my_FIR_filter_firBlock_left_add_221_carry[11]), .YC(my_FIR_filter_firBlock_left_add_221_carry[12]), .YS(my_FIR_filter_firBlock_left_N44));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_12 ( .A(n442),  .B(my_FIR_filter_firBlock_left_multProducts[45]),  .C(my_FIR_filter_firBlock_left_add_221_carry[12]), .YC(my_FIR_filter_firBlock_left_add_221_carry[13]), .YS(my_FIR_filter_firBlock_left_N45));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_13 ( .A(n443),  .B(my_FIR_filter_firBlock_left_multProducts[46]),  .C(my_FIR_filter_firBlock_left_add_221_carry[13]), .YC(my_FIR_filter_firBlock_left_add_221_carry[14]), .YS(my_FIR_filter_firBlock_left_N46));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_14 ( .A(n444),  .B(my_FIR_filter_firBlock_left_multProducts[47]),  .C(my_FIR_filter_firBlock_left_add_221_carry[14]), .YC(my_FIR_filter_firBlock_left_add_221_carry[15]), .YS(my_FIR_filter_firBlock_left_N47));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_15 ( .A(n445),  .B(my_FIR_filter_firBlock_left_multProducts[48]),  .C(my_FIR_filter_firBlock_left_add_221_carry[15]), .YC(my_FIR_filter_firBlock_left_add_221_carry[16]), .YS(my_FIR_filter_firBlock_left_N48));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_16 ( .A(n446),  .B(my_FIR_filter_firBlock_left_multProducts[49]),  .C(my_FIR_filter_firBlock_left_add_221_carry[16]), .YC(my_FIR_filter_firBlock_left_add_221_carry[17]), .YS(my_FIR_filter_firBlock_left_N49));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_17 ( .A(n447),  .B(my_FIR_filter_firBlock_left_multProducts[50]),  .C(my_FIR_filter_firBlock_left_add_221_carry[17]), .YC(my_FIR_filter_firBlock_left_add_221_carry[18]), .YS(my_FIR_filter_firBlock_left_N50));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_18 ( .A(n448),  .B(my_FIR_filter_firBlock_left_multProducts[51]),  .C(my_FIR_filter_firBlock_left_add_221_carry[18]), .YC(my_FIR_filter_firBlock_left_add_221_carry[19]), .YS(my_FIR_filter_firBlock_left_N51));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_19 ( .A(n449),  .B(my_FIR_filter_firBlock_left_multProducts[52]),  .C(my_FIR_filter_firBlock_left_add_221_carry[19]), .YC(my_FIR_filter_firBlock_left_add_221_carry[20]), .YS(my_FIR_filter_firBlock_left_N52));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_20 ( .A(n450),  .B(my_FIR_filter_firBlock_left_multProducts[53]),  .C(my_FIR_filter_firBlock_left_add_221_carry[20]), .YC(my_FIR_filter_firBlock_left_add_221_carry[21]), .YS(my_FIR_filter_firBlock_left_N53));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_21 ( .A(n451),  .B(my_FIR_filter_firBlock_left_multProducts[54]),  .C(my_FIR_filter_firBlock_left_add_221_carry[21]), .YC(my_FIR_filter_firBlock_left_add_221_carry[22]), .YS(my_FIR_filter_firBlock_left_N54));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_22 ( .A(n452),  .B(my_FIR_filter_firBlock_left_multProducts[55]),  .C(my_FIR_filter_firBlock_left_add_221_carry[22]), .YC(my_FIR_filter_firBlock_left_add_221_carry[23]), .YS(my_FIR_filter_firBlock_left_N55));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_23 ( .A(n453),  .B(my_FIR_filter_firBlock_left_multProducts[56]),  .C(my_FIR_filter_firBlock_left_add_221_carry[23]), .YC(my_FIR_filter_firBlock_left_add_221_carry[24]), .YS(my_FIR_filter_firBlock_left_N56));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_24 ( .A(n454),  .B(my_FIR_filter_firBlock_left_multProducts[57]),  .C(my_FIR_filter_firBlock_left_add_221_carry[24]), .YC(my_FIR_filter_firBlock_left_add_221_carry[25]), .YS(my_FIR_filter_firBlock_left_N57));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_25 ( .A(n455),  .B(my_FIR_filter_firBlock_left_multProducts[58]),  .C(my_FIR_filter_firBlock_left_add_221_carry[25]), .YC(my_FIR_filter_firBlock_left_add_221_carry[26]), .YS(my_FIR_filter_firBlock_left_N58));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_26 ( .A(n456),  .B(my_FIR_filter_firBlock_left_multProducts[59]),  .C(my_FIR_filter_firBlock_left_add_221_carry[26]), .YC(my_FIR_filter_firBlock_left_add_221_carry[27]), .YS(my_FIR_filter_firBlock_left_N59));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_27 ( .A(n457),  .B(my_FIR_filter_firBlock_left_multProducts[60]),  .C(my_FIR_filter_firBlock_left_add_221_carry[27]), .YC(my_FIR_filter_firBlock_left_add_221_carry[28]), .YS(my_FIR_filter_firBlock_left_N60));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_28 ( .A(n458),  .B(my_FIR_filter_firBlock_left_multProducts[61]),  .C(my_FIR_filter_firBlock_left_add_221_carry[28]), .YC(my_FIR_filter_firBlock_left_add_221_carry[29]), .YS(my_FIR_filter_firBlock_left_N61));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_29 ( .A(n459),  .B(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[35]),  .C(my_FIR_filter_firBlock_left_add_221_carry[29]), .YC(my_FIR_filter_firBlock_left_add_221_carry[30]), .YS(my_FIR_filter_firBlock_left_N62));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_30 ( .A(n121),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_221_carry[30]), .YC(my_FIR_filter_firBlock_left_add_221_carry[31]), .YS(my_FIR_filter_firBlock_left_N63));
   FAX1 my_FIR_filter_firBlock_left_add_221_U1_31 ( .A(n122),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_221_carry[31]), .YS(my_FIR_filter_firBlock_left_N64));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_1 ( .A(n297),  .B(my_FIR_filter_firBlock_left_multProducts[33]),  .C(n520), .YC(my_FIR_filter_firBlock_left_add_222_carry[2]), .YS(my_FIR_filter_firBlock_left_N66));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_2 ( .A(n246),  .B(my_FIR_filter_firBlock_left_multProducts[34]),  .C(my_FIR_filter_firBlock_left_add_222_carry[2]), .YC(my_FIR_filter_firBlock_left_add_222_carry[3]), .YS(my_FIR_filter_firBlock_left_N67));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_3 ( .A(n247),  .B(my_FIR_filter_firBlock_left_multProducts[35]),  .C(my_FIR_filter_firBlock_left_add_222_carry[3]), .YC(my_FIR_filter_firBlock_left_add_222_carry[4]), .YS(my_FIR_filter_firBlock_left_N68));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_4 ( .A(n248),  .B(my_FIR_filter_firBlock_left_multProducts[36]),  .C(my_FIR_filter_firBlock_left_add_222_carry[4]), .YC(my_FIR_filter_firBlock_left_add_222_carry[5]), .YS(my_FIR_filter_firBlock_left_N69));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_5 ( .A(n249),  .B(my_FIR_filter_firBlock_left_multProducts[37]),  .C(my_FIR_filter_firBlock_left_add_222_carry[5]), .YC(my_FIR_filter_firBlock_left_add_222_carry[6]), .YS(my_FIR_filter_firBlock_left_N70));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_6 ( .A(n250),  .B(my_FIR_filter_firBlock_left_multProducts[38]),  .C(my_FIR_filter_firBlock_left_add_222_carry[6]), .YC(my_FIR_filter_firBlock_left_add_222_carry[7]), .YS(my_FIR_filter_firBlock_left_N71));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_7 ( .A(n251),  .B(my_FIR_filter_firBlock_left_multProducts[39]),  .C(my_FIR_filter_firBlock_left_add_222_carry[7]), .YC(my_FIR_filter_firBlock_left_add_222_carry[8]), .YS(my_FIR_filter_firBlock_left_N72));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_8 ( .A(n252),  .B(my_FIR_filter_firBlock_left_multProducts[40]),  .C(my_FIR_filter_firBlock_left_add_222_carry[8]), .YC(my_FIR_filter_firBlock_left_add_222_carry[9]), .YS(my_FIR_filter_firBlock_left_N73));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_9 ( .A(n253),  .B(my_FIR_filter_firBlock_left_multProducts[41]),  .C(my_FIR_filter_firBlock_left_add_222_carry[9]), .YC(my_FIR_filter_firBlock_left_add_222_carry[10]), .YS(my_FIR_filter_firBlock_left_N74));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_10 ( .A(n254),  .B(my_FIR_filter_firBlock_left_multProducts[42]),  .C(my_FIR_filter_firBlock_left_add_222_carry[10]), .YC(my_FIR_filter_firBlock_left_add_222_carry[11]), .YS(my_FIR_filter_firBlock_left_N75));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_11 ( .A(n255),  .B(my_FIR_filter_firBlock_left_multProducts[43]),  .C(my_FIR_filter_firBlock_left_add_222_carry[11]), .YC(my_FIR_filter_firBlock_left_add_222_carry[12]), .YS(my_FIR_filter_firBlock_left_N76));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_12 ( .A(n256),  .B(my_FIR_filter_firBlock_left_multProducts[44]),  .C(my_FIR_filter_firBlock_left_add_222_carry[12]), .YC(my_FIR_filter_firBlock_left_add_222_carry[13]), .YS(my_FIR_filter_firBlock_left_N77));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_13 ( .A(n257),  .B(my_FIR_filter_firBlock_left_multProducts[45]),  .C(my_FIR_filter_firBlock_left_add_222_carry[13]), .YC(my_FIR_filter_firBlock_left_add_222_carry[14]), .YS(my_FIR_filter_firBlock_left_N78));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_14 ( .A(n258),  .B(my_FIR_filter_firBlock_left_multProducts[46]),  .C(my_FIR_filter_firBlock_left_add_222_carry[14]), .YC(my_FIR_filter_firBlock_left_add_222_carry[15]), .YS(my_FIR_filter_firBlock_left_N79));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_15 ( .A(n259),  .B(my_FIR_filter_firBlock_left_multProducts[47]),  .C(my_FIR_filter_firBlock_left_add_222_carry[15]), .YC(my_FIR_filter_firBlock_left_add_222_carry[16]), .YS(my_FIR_filter_firBlock_left_N80));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_16 ( .A(n260),  .B(my_FIR_filter_firBlock_left_multProducts[48]),  .C(my_FIR_filter_firBlock_left_add_222_carry[16]), .YC(my_FIR_filter_firBlock_left_add_222_carry[17]), .YS(my_FIR_filter_firBlock_left_N81));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_17 ( .A(n261),  .B(my_FIR_filter_firBlock_left_multProducts[49]),  .C(my_FIR_filter_firBlock_left_add_222_carry[17]), .YC(my_FIR_filter_firBlock_left_add_222_carry[18]), .YS(my_FIR_filter_firBlock_left_N82));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_18 ( .A(n262),  .B(my_FIR_filter_firBlock_left_multProducts[50]),  .C(my_FIR_filter_firBlock_left_add_222_carry[18]), .YC(my_FIR_filter_firBlock_left_add_222_carry[19]), .YS(my_FIR_filter_firBlock_left_N83));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_19 ( .A(n263),  .B(my_FIR_filter_firBlock_left_multProducts[51]),  .C(my_FIR_filter_firBlock_left_add_222_carry[19]), .YC(my_FIR_filter_firBlock_left_add_222_carry[20]), .YS(my_FIR_filter_firBlock_left_N84));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_20 ( .A(n264),  .B(my_FIR_filter_firBlock_left_multProducts[52]),  .C(my_FIR_filter_firBlock_left_add_222_carry[20]), .YC(my_FIR_filter_firBlock_left_add_222_carry[21]), .YS(my_FIR_filter_firBlock_left_N85));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_21 ( .A(n265),  .B(my_FIR_filter_firBlock_left_multProducts[53]),  .C(my_FIR_filter_firBlock_left_add_222_carry[21]), .YC(my_FIR_filter_firBlock_left_add_222_carry[22]), .YS(my_FIR_filter_firBlock_left_N86));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_22 ( .A(n266),  .B(my_FIR_filter_firBlock_left_multProducts[54]),  .C(my_FIR_filter_firBlock_left_add_222_carry[22]), .YC(my_FIR_filter_firBlock_left_add_222_carry[23]), .YS(my_FIR_filter_firBlock_left_N87));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_23 ( .A(n267),  .B(my_FIR_filter_firBlock_left_multProducts[55]),  .C(my_FIR_filter_firBlock_left_add_222_carry[23]), .YC(my_FIR_filter_firBlock_left_add_222_carry[24]), .YS(my_FIR_filter_firBlock_left_N88));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_24 ( .A(n268),  .B(my_FIR_filter_firBlock_left_multProducts[56]),  .C(my_FIR_filter_firBlock_left_add_222_carry[24]), .YC(my_FIR_filter_firBlock_left_add_222_carry[25]), .YS(my_FIR_filter_firBlock_left_N89));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_25 ( .A(n269),  .B(my_FIR_filter_firBlock_left_multProducts[57]),  .C(my_FIR_filter_firBlock_left_add_222_carry[25]), .YC(my_FIR_filter_firBlock_left_add_222_carry[26]), .YS(my_FIR_filter_firBlock_left_N90));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_26 ( .A(n270),  .B(my_FIR_filter_firBlock_left_multProducts[58]),  .C(my_FIR_filter_firBlock_left_add_222_carry[26]), .YC(my_FIR_filter_firBlock_left_add_222_carry[27]), .YS(my_FIR_filter_firBlock_left_N91));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_27 ( .A(n271),  .B(my_FIR_filter_firBlock_left_multProducts[59]),  .C(my_FIR_filter_firBlock_left_add_222_carry[27]), .YC(my_FIR_filter_firBlock_left_add_222_carry[28]), .YS(my_FIR_filter_firBlock_left_N92));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_28 ( .A(n272),  .B(my_FIR_filter_firBlock_left_multProducts[60]),  .C(my_FIR_filter_firBlock_left_add_222_carry[28]), .YC(my_FIR_filter_firBlock_left_add_222_carry[29]), .YS(my_FIR_filter_firBlock_left_N93));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_29 ( .A(n273),  .B(my_FIR_filter_firBlock_left_multProducts[61]),  .C(my_FIR_filter_firBlock_left_add_222_carry[29]), .YC(my_FIR_filter_firBlock_left_add_222_carry[30]), .YS(my_FIR_filter_firBlock_left_N94));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_30 ( .A(n274),  .B(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[35]),  .C(my_FIR_filter_firBlock_left_add_222_carry[30]), .YC(my_FIR_filter_firBlock_left_add_222_carry[31]), .YS(my_FIR_filter_firBlock_left_N95));
   FAX1 my_FIR_filter_firBlock_left_add_222_U1_31 ( .A(n275),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_222_carry[31]), .YS(my_FIR_filter_firBlock_left_N96));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_1 ( .A(n466),  .B(my_FIR_filter_firBlock_left_multProducts[1]),  .C(n521), .YC(my_FIR_filter_firBlock_left_add_223_carry[2]), .YS(my_FIR_filter_firBlock_left_N98));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_2 ( .A(n403),  .B(my_FIR_filter_firBlock_left_multProducts[2]),  .C(my_FIR_filter_firBlock_left_add_223_carry[2]), .YC(my_FIR_filter_firBlock_left_add_223_carry[3]), .YS(my_FIR_filter_firBlock_left_N99));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_3 ( .A(n404),  .B(my_FIR_filter_firBlock_left_multProducts[3]),  .C(my_FIR_filter_firBlock_left_add_223_carry[3]), .YC(my_FIR_filter_firBlock_left_add_223_carry[4]), .YS(my_FIR_filter_firBlock_left_N100));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_4 ( .A(n405),  .B(my_FIR_filter_firBlock_left_multProducts[4]),  .C(my_FIR_filter_firBlock_left_add_223_carry[4]), .YC(my_FIR_filter_firBlock_left_add_223_carry[5]), .YS(my_FIR_filter_firBlock_left_N101));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_5 ( .A(n406),  .B(my_FIR_filter_firBlock_left_multProducts[5]),  .C(my_FIR_filter_firBlock_left_add_223_carry[5]), .YC(my_FIR_filter_firBlock_left_add_223_carry[6]), .YS(my_FIR_filter_firBlock_left_N102));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_6 ( .A(n407),  .B(my_FIR_filter_firBlock_left_multProducts[6]),  .C(my_FIR_filter_firBlock_left_add_223_carry[6]), .YC(my_FIR_filter_firBlock_left_add_223_carry[7]), .YS(my_FIR_filter_firBlock_left_N103));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_7 ( .A(n408),  .B(my_FIR_filter_firBlock_left_multProducts[7]),  .C(my_FIR_filter_firBlock_left_add_223_carry[7]), .YC(my_FIR_filter_firBlock_left_add_223_carry[8]), .YS(my_FIR_filter_firBlock_left_N104));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_8 ( .A(n409),  .B(my_FIR_filter_firBlock_left_multProducts[8]),  .C(my_FIR_filter_firBlock_left_add_223_carry[8]), .YC(my_FIR_filter_firBlock_left_add_223_carry[9]), .YS(my_FIR_filter_firBlock_left_N105));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_9 ( .A(n410),  .B(my_FIR_filter_firBlock_left_multProducts[9]),  .C(my_FIR_filter_firBlock_left_add_223_carry[9]), .YC(my_FIR_filter_firBlock_left_add_223_carry[10]), .YS(my_FIR_filter_firBlock_left_N106));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_10 ( .A(n411),  .B(my_FIR_filter_firBlock_left_multProducts[10]),  .C(my_FIR_filter_firBlock_left_add_223_carry[10]), .YC(my_FIR_filter_firBlock_left_add_223_carry[11]), .YS(my_FIR_filter_firBlock_left_N107));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_11 ( .A(n412),  .B(my_FIR_filter_firBlock_left_multProducts[11]),  .C(my_FIR_filter_firBlock_left_add_223_carry[11]), .YC(my_FIR_filter_firBlock_left_add_223_carry[12]), .YS(my_FIR_filter_firBlock_left_N108));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_12 ( .A(n413),  .B(my_FIR_filter_firBlock_left_multProducts[12]),  .C(my_FIR_filter_firBlock_left_add_223_carry[12]), .YC(my_FIR_filter_firBlock_left_add_223_carry[13]), .YS(my_FIR_filter_firBlock_left_N109));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_13 ( .A(n414),  .B(my_FIR_filter_firBlock_left_multProducts[13]),  .C(my_FIR_filter_firBlock_left_add_223_carry[13]), .YC(my_FIR_filter_firBlock_left_add_223_carry[14]), .YS(my_FIR_filter_firBlock_left_N110));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_14 ( .A(n415),  .B(my_FIR_filter_firBlock_left_multProducts[14]),  .C(my_FIR_filter_firBlock_left_add_223_carry[14]), .YC(my_FIR_filter_firBlock_left_add_223_carry[15]), .YS(my_FIR_filter_firBlock_left_N111));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_15 ( .A(n416),  .B(my_FIR_filter_firBlock_left_multProducts[15]),  .C(my_FIR_filter_firBlock_left_add_223_carry[15]), .YC(my_FIR_filter_firBlock_left_add_223_carry[16]), .YS(my_FIR_filter_firBlock_left_N112));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_16 ( .A(n417),  .B(my_FIR_filter_firBlock_left_multProducts[16]),  .C(my_FIR_filter_firBlock_left_add_223_carry[16]), .YC(my_FIR_filter_firBlock_left_add_223_carry[17]), .YS(my_FIR_filter_firBlock_left_N113));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_17 ( .A(n418),  .B(my_FIR_filter_firBlock_left_multProducts[17]),  .C(my_FIR_filter_firBlock_left_add_223_carry[17]), .YC(my_FIR_filter_firBlock_left_add_223_carry[18]), .YS(my_FIR_filter_firBlock_left_N114));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_18 ( .A(n419),  .B(my_FIR_filter_firBlock_left_multProducts[18]),  .C(my_FIR_filter_firBlock_left_add_223_carry[18]), .YC(my_FIR_filter_firBlock_left_add_223_carry[19]), .YS(my_FIR_filter_firBlock_left_N115));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_19 ( .A(n420),  .B(my_FIR_filter_firBlock_left_multProducts[19]),  .C(my_FIR_filter_firBlock_left_add_223_carry[19]), .YC(my_FIR_filter_firBlock_left_add_223_carry[20]), .YS(my_FIR_filter_firBlock_left_N116));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_20 ( .A(n421),  .B(my_FIR_filter_firBlock_left_multProducts[20]),  .C(my_FIR_filter_firBlock_left_add_223_carry[20]), .YC(my_FIR_filter_firBlock_left_add_223_carry[21]), .YS(my_FIR_filter_firBlock_left_N117));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_21 ( .A(n422),  .B(my_FIR_filter_firBlock_left_multProducts[21]),  .C(my_FIR_filter_firBlock_left_add_223_carry[21]), .YC(my_FIR_filter_firBlock_left_add_223_carry[22]), .YS(my_FIR_filter_firBlock_left_N118));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_22 ( .A(n423),  .B(my_FIR_filter_firBlock_left_multProducts[22]),  .C(my_FIR_filter_firBlock_left_add_223_carry[22]), .YC(my_FIR_filter_firBlock_left_add_223_carry[23]), .YS(my_FIR_filter_firBlock_left_N119));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_23 ( .A(n424),  .B(my_FIR_filter_firBlock_left_multProducts[23]),  .C(my_FIR_filter_firBlock_left_add_223_carry[23]), .YC(my_FIR_filter_firBlock_left_add_223_carry[24]), .YS(my_FIR_filter_firBlock_left_N120));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_24 ( .A(n425),  .B(my_FIR_filter_firBlock_left_multProducts[24]),  .C(my_FIR_filter_firBlock_left_add_223_carry[24]), .YC(my_FIR_filter_firBlock_left_add_223_carry[25]), .YS(my_FIR_filter_firBlock_left_N121));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_25 ( .A(n426),  .B(my_FIR_filter_firBlock_left_multProducts[25]),  .C(my_FIR_filter_firBlock_left_add_223_carry[25]), .YC(my_FIR_filter_firBlock_left_add_223_carry[26]), .YS(my_FIR_filter_firBlock_left_N122));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_26 ( .A(n427),  .B(my_FIR_filter_firBlock_left_multProducts[26]),  .C(my_FIR_filter_firBlock_left_add_223_carry[26]), .YC(my_FIR_filter_firBlock_left_add_223_carry[27]), .YS(my_FIR_filter_firBlock_left_N123));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_27 ( .A(n428),  .B(my_FIR_filter_firBlock_left_multProducts[27]),  .C(my_FIR_filter_firBlock_left_add_223_carry[27]), .YC(my_FIR_filter_firBlock_left_add_223_carry[28]), .YS(my_FIR_filter_firBlock_left_N124));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_28 ( .A(n429),  .B(my_FIR_filter_firBlock_left_multProducts[28]),  .C(my_FIR_filter_firBlock_left_add_223_carry[28]), .YC(my_FIR_filter_firBlock_left_add_223_carry[29]), .YS(my_FIR_filter_firBlock_left_N125));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_29 ( .A(n430),  .B(my_FIR_filter_firBlock_left_multProducts[29]),  .C(my_FIR_filter_firBlock_left_add_223_carry[29]), .YC(my_FIR_filter_firBlock_left_add_223_carry[30]), .YS(my_FIR_filter_firBlock_left_N126));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_30 ( .A(n431),  .B(my_FIR_filter_firBlock_left_multProducts[30]),  .C(my_FIR_filter_firBlock_left_add_223_carry[30]), .YC(my_FIR_filter_firBlock_left_add_223_carry[31]), .YS(my_FIR_filter_firBlock_left_N127));
   FAX1 my_FIR_filter_firBlock_left_add_223_U1_31 ( .A(n120),  .B(my_FIR_filter_firBlock_left_multProducts[31]),  .C(my_FIR_filter_firBlock_left_add_223_carry[31]), .YS(my_FIR_filter_firBlock_left_N128));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_1 ( .A(n296),  .B(my_FIR_filter_firBlock_left_multProducts[1]),  .C(n522), .YC(my_FIR_filter_firBlock_left_add_224_carry[2]), .YS(my_FIR_filter_firBlock_left_N130));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_2 ( .A(n217),  .B(my_FIR_filter_firBlock_left_multProducts[2]),  .C(my_FIR_filter_firBlock_left_add_224_carry[2]), .YC(my_FIR_filter_firBlock_left_add_224_carry[3]), .YS(my_FIR_filter_firBlock_left_N131));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_3 ( .A(n218),  .B(my_FIR_filter_firBlock_left_multProducts[3]),  .C(my_FIR_filter_firBlock_left_add_224_carry[3]), .YC(my_FIR_filter_firBlock_left_add_224_carry[4]), .YS(my_FIR_filter_firBlock_left_N132));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_4 ( .A(n219),  .B(my_FIR_filter_firBlock_left_multProducts[4]),  .C(my_FIR_filter_firBlock_left_add_224_carry[4]), .YC(my_FIR_filter_firBlock_left_add_224_carry[5]), .YS(my_FIR_filter_firBlock_left_N133));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_5 ( .A(n220),  .B(my_FIR_filter_firBlock_left_multProducts[5]),  .C(my_FIR_filter_firBlock_left_add_224_carry[5]), .YC(my_FIR_filter_firBlock_left_add_224_carry[6]), .YS(my_FIR_filter_firBlock_left_N134));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_6 ( .A(n221),  .B(my_FIR_filter_firBlock_left_multProducts[6]),  .C(my_FIR_filter_firBlock_left_add_224_carry[6]), .YC(my_FIR_filter_firBlock_left_add_224_carry[7]), .YS(my_FIR_filter_firBlock_left_N135));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_7 ( .A(n222),  .B(my_FIR_filter_firBlock_left_multProducts[7]),  .C(my_FIR_filter_firBlock_left_add_224_carry[7]), .YC(my_FIR_filter_firBlock_left_add_224_carry[8]), .YS(my_FIR_filter_firBlock_left_N136));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_8 ( .A(n223),  .B(my_FIR_filter_firBlock_left_multProducts[8]),  .C(my_FIR_filter_firBlock_left_add_224_carry[8]), .YC(my_FIR_filter_firBlock_left_add_224_carry[9]), .YS(my_FIR_filter_firBlock_left_N137));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_9 ( .A(n224),  .B(my_FIR_filter_firBlock_left_multProducts[9]),  .C(my_FIR_filter_firBlock_left_add_224_carry[9]), .YC(my_FIR_filter_firBlock_left_add_224_carry[10]), .YS(my_FIR_filter_firBlock_left_N138));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_10 ( .A(n225),  .B(my_FIR_filter_firBlock_left_multProducts[10]),  .C(my_FIR_filter_firBlock_left_add_224_carry[10]), .YC(my_FIR_filter_firBlock_left_add_224_carry[11]), .YS(my_FIR_filter_firBlock_left_N139));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_11 ( .A(n226),  .B(my_FIR_filter_firBlock_left_multProducts[11]),  .C(my_FIR_filter_firBlock_left_add_224_carry[11]), .YC(my_FIR_filter_firBlock_left_add_224_carry[12]), .YS(my_FIR_filter_firBlock_left_N140));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_12 ( .A(n227),  .B(my_FIR_filter_firBlock_left_multProducts[12]),  .C(my_FIR_filter_firBlock_left_add_224_carry[12]), .YC(my_FIR_filter_firBlock_left_add_224_carry[13]), .YS(my_FIR_filter_firBlock_left_N141));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_13 ( .A(n228),  .B(my_FIR_filter_firBlock_left_multProducts[13]),  .C(my_FIR_filter_firBlock_left_add_224_carry[13]), .YC(my_FIR_filter_firBlock_left_add_224_carry[14]), .YS(my_FIR_filter_firBlock_left_N142));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_14 ( .A(n229),  .B(my_FIR_filter_firBlock_left_multProducts[14]),  .C(my_FIR_filter_firBlock_left_add_224_carry[14]), .YC(my_FIR_filter_firBlock_left_add_224_carry[15]), .YS(my_FIR_filter_firBlock_left_N143));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_15 ( .A(n230),  .B(my_FIR_filter_firBlock_left_multProducts[15]),  .C(my_FIR_filter_firBlock_left_add_224_carry[15]), .YC(my_FIR_filter_firBlock_left_add_224_carry[16]), .YS(my_FIR_filter_firBlock_left_N144));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_16 ( .A(n231),  .B(my_FIR_filter_firBlock_left_multProducts[16]),  .C(my_FIR_filter_firBlock_left_add_224_carry[16]), .YC(my_FIR_filter_firBlock_left_add_224_carry[17]), .YS(my_FIR_filter_firBlock_left_N145));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_17 ( .A(n232),  .B(my_FIR_filter_firBlock_left_multProducts[17]),  .C(my_FIR_filter_firBlock_left_add_224_carry[17]), .YC(my_FIR_filter_firBlock_left_add_224_carry[18]), .YS(my_FIR_filter_firBlock_left_N146));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_18 ( .A(n233),  .B(my_FIR_filter_firBlock_left_multProducts[18]),  .C(my_FIR_filter_firBlock_left_add_224_carry[18]), .YC(my_FIR_filter_firBlock_left_add_224_carry[19]), .YS(my_FIR_filter_firBlock_left_N147));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_19 ( .A(n234),  .B(my_FIR_filter_firBlock_left_multProducts[19]),  .C(my_FIR_filter_firBlock_left_add_224_carry[19]), .YC(my_FIR_filter_firBlock_left_add_224_carry[20]), .YS(my_FIR_filter_firBlock_left_N148));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_20 ( .A(n235),  .B(my_FIR_filter_firBlock_left_multProducts[20]),  .C(my_FIR_filter_firBlock_left_add_224_carry[20]), .YC(my_FIR_filter_firBlock_left_add_224_carry[21]), .YS(my_FIR_filter_firBlock_left_N149));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_21 ( .A(n236),  .B(my_FIR_filter_firBlock_left_multProducts[21]),  .C(my_FIR_filter_firBlock_left_add_224_carry[21]), .YC(my_FIR_filter_firBlock_left_add_224_carry[22]), .YS(my_FIR_filter_firBlock_left_N150));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_22 ( .A(n237),  .B(my_FIR_filter_firBlock_left_multProducts[22]),  .C(my_FIR_filter_firBlock_left_add_224_carry[22]), .YC(my_FIR_filter_firBlock_left_add_224_carry[23]), .YS(my_FIR_filter_firBlock_left_N151));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_23 ( .A(n238),  .B(my_FIR_filter_firBlock_left_multProducts[23]),  .C(my_FIR_filter_firBlock_left_add_224_carry[23]), .YC(my_FIR_filter_firBlock_left_add_224_carry[24]), .YS(my_FIR_filter_firBlock_left_N152));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_24 ( .A(n239),  .B(my_FIR_filter_firBlock_left_multProducts[24]),  .C(my_FIR_filter_firBlock_left_add_224_carry[24]), .YC(my_FIR_filter_firBlock_left_add_224_carry[25]), .YS(my_FIR_filter_firBlock_left_N153));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_25 ( .A(n240),  .B(my_FIR_filter_firBlock_left_multProducts[25]),  .C(my_FIR_filter_firBlock_left_add_224_carry[25]), .YC(my_FIR_filter_firBlock_left_add_224_carry[26]), .YS(my_FIR_filter_firBlock_left_N154));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_26 ( .A(n241),  .B(my_FIR_filter_firBlock_left_multProducts[26]),  .C(my_FIR_filter_firBlock_left_add_224_carry[26]), .YC(my_FIR_filter_firBlock_left_add_224_carry[27]), .YS(my_FIR_filter_firBlock_left_N155));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_27 ( .A(n242),  .B(my_FIR_filter_firBlock_left_multProducts[27]),  .C(my_FIR_filter_firBlock_left_add_224_carry[27]), .YC(my_FIR_filter_firBlock_left_add_224_carry[28]), .YS(my_FIR_filter_firBlock_left_N156));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_28 ( .A(n243),  .B(my_FIR_filter_firBlock_left_multProducts[28]),  .C(my_FIR_filter_firBlock_left_add_224_carry[28]), .YC(my_FIR_filter_firBlock_left_add_224_carry[29]), .YS(my_FIR_filter_firBlock_left_N157));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_29 ( .A(n244),  .B(my_FIR_filter_firBlock_left_multProducts[29]),  .C(my_FIR_filter_firBlock_left_add_224_carry[29]), .YC(my_FIR_filter_firBlock_left_add_224_carry[30]), .YS(my_FIR_filter_firBlock_left_N158));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_30 ( .A(n245),  .B(my_FIR_filter_firBlock_left_multProducts[30]),  .C(my_FIR_filter_firBlock_left_add_224_carry[30]), .YC(my_FIR_filter_firBlock_left_add_224_carry[31]), .YS(my_FIR_filter_firBlock_left_N159));
   FAX1 my_FIR_filter_firBlock_left_add_224_U1_31 ( .A(n402),  .B(my_FIR_filter_firBlock_left_multProducts[31]),  .C(my_FIR_filter_firBlock_left_add_224_carry[31]), .YS(my_FIR_filter_firBlock_left_N160));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_1 ( .A(n465),  .B(my_FIR_filter_firBlock_left_multProducts[33]),  .C(n523), .YC(my_FIR_filter_firBlock_left_add_225_carry[2]), .YS(my_FIR_filter_firBlock_left_N162));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_2 ( .A(n373),  .B(my_FIR_filter_firBlock_left_multProducts[34]),  .C(my_FIR_filter_firBlock_left_add_225_carry[2]), .YC(my_FIR_filter_firBlock_left_add_225_carry[3]), .YS(my_FIR_filter_firBlock_left_N163));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_3 ( .A(n374),  .B(my_FIR_filter_firBlock_left_multProducts[35]),  .C(my_FIR_filter_firBlock_left_add_225_carry[3]), .YC(my_FIR_filter_firBlock_left_add_225_carry[4]), .YS(my_FIR_filter_firBlock_left_N164));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_4 ( .A(n375),  .B(my_FIR_filter_firBlock_left_multProducts[36]),  .C(my_FIR_filter_firBlock_left_add_225_carry[4]), .YC(my_FIR_filter_firBlock_left_add_225_carry[5]), .YS(my_FIR_filter_firBlock_left_N165));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_5 ( .A(n376),  .B(my_FIR_filter_firBlock_left_multProducts[37]),  .C(my_FIR_filter_firBlock_left_add_225_carry[5]), .YC(my_FIR_filter_firBlock_left_add_225_carry[6]), .YS(my_FIR_filter_firBlock_left_N166));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_6 ( .A(n377),  .B(my_FIR_filter_firBlock_left_multProducts[38]),  .C(my_FIR_filter_firBlock_left_add_225_carry[6]), .YC(my_FIR_filter_firBlock_left_add_225_carry[7]), .YS(my_FIR_filter_firBlock_left_N167));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_7 ( .A(n378),  .B(my_FIR_filter_firBlock_left_multProducts[39]),  .C(my_FIR_filter_firBlock_left_add_225_carry[7]), .YC(my_FIR_filter_firBlock_left_add_225_carry[8]), .YS(my_FIR_filter_firBlock_left_N168));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_8 ( .A(n379),  .B(my_FIR_filter_firBlock_left_multProducts[40]),  .C(my_FIR_filter_firBlock_left_add_225_carry[8]), .YC(my_FIR_filter_firBlock_left_add_225_carry[9]), .YS(my_FIR_filter_firBlock_left_N169));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_9 ( .A(n380),  .B(my_FIR_filter_firBlock_left_multProducts[41]),  .C(my_FIR_filter_firBlock_left_add_225_carry[9]), .YC(my_FIR_filter_firBlock_left_add_225_carry[10]), .YS(my_FIR_filter_firBlock_left_N170));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_10 ( .A(n381),  .B(my_FIR_filter_firBlock_left_multProducts[42]),  .C(my_FIR_filter_firBlock_left_add_225_carry[10]), .YC(my_FIR_filter_firBlock_left_add_225_carry[11]), .YS(my_FIR_filter_firBlock_left_N171));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_11 ( .A(n382),  .B(my_FIR_filter_firBlock_left_multProducts[43]),  .C(my_FIR_filter_firBlock_left_add_225_carry[11]), .YC(my_FIR_filter_firBlock_left_add_225_carry[12]), .YS(my_FIR_filter_firBlock_left_N172));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_12 ( .A(n383),  .B(my_FIR_filter_firBlock_left_multProducts[44]),  .C(my_FIR_filter_firBlock_left_add_225_carry[12]), .YC(my_FIR_filter_firBlock_left_add_225_carry[13]), .YS(my_FIR_filter_firBlock_left_N173));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_13 ( .A(n384),  .B(my_FIR_filter_firBlock_left_multProducts[45]),  .C(my_FIR_filter_firBlock_left_add_225_carry[13]), .YC(my_FIR_filter_firBlock_left_add_225_carry[14]), .YS(my_FIR_filter_firBlock_left_N174));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_14 ( .A(n385),  .B(my_FIR_filter_firBlock_left_multProducts[46]),  .C(my_FIR_filter_firBlock_left_add_225_carry[14]), .YC(my_FIR_filter_firBlock_left_add_225_carry[15]), .YS(my_FIR_filter_firBlock_left_N175));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_15 ( .A(n386),  .B(my_FIR_filter_firBlock_left_multProducts[47]),  .C(my_FIR_filter_firBlock_left_add_225_carry[15]), .YC(my_FIR_filter_firBlock_left_add_225_carry[16]), .YS(my_FIR_filter_firBlock_left_N176));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_16 ( .A(n387),  .B(my_FIR_filter_firBlock_left_multProducts[48]),  .C(my_FIR_filter_firBlock_left_add_225_carry[16]), .YC(my_FIR_filter_firBlock_left_add_225_carry[17]), .YS(my_FIR_filter_firBlock_left_N177));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_17 ( .A(n388),  .B(my_FIR_filter_firBlock_left_multProducts[49]),  .C(my_FIR_filter_firBlock_left_add_225_carry[17]), .YC(my_FIR_filter_firBlock_left_add_225_carry[18]), .YS(my_FIR_filter_firBlock_left_N178));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_18 ( .A(n389),  .B(my_FIR_filter_firBlock_left_multProducts[50]),  .C(my_FIR_filter_firBlock_left_add_225_carry[18]), .YC(my_FIR_filter_firBlock_left_add_225_carry[19]), .YS(my_FIR_filter_firBlock_left_N179));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_19 ( .A(n390),  .B(my_FIR_filter_firBlock_left_multProducts[51]),  .C(my_FIR_filter_firBlock_left_add_225_carry[19]), .YC(my_FIR_filter_firBlock_left_add_225_carry[20]), .YS(my_FIR_filter_firBlock_left_N180));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_20 ( .A(n391),  .B(my_FIR_filter_firBlock_left_multProducts[52]),  .C(my_FIR_filter_firBlock_left_add_225_carry[20]), .YC(my_FIR_filter_firBlock_left_add_225_carry[21]), .YS(my_FIR_filter_firBlock_left_N181));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_21 ( .A(n392),  .B(my_FIR_filter_firBlock_left_multProducts[53]),  .C(my_FIR_filter_firBlock_left_add_225_carry[21]), .YC(my_FIR_filter_firBlock_left_add_225_carry[22]), .YS(my_FIR_filter_firBlock_left_N182));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_22 ( .A(n393),  .B(my_FIR_filter_firBlock_left_multProducts[54]),  .C(my_FIR_filter_firBlock_left_add_225_carry[22]), .YC(my_FIR_filter_firBlock_left_add_225_carry[23]), .YS(my_FIR_filter_firBlock_left_N183));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_23 ( .A(n394),  .B(my_FIR_filter_firBlock_left_multProducts[55]),  .C(my_FIR_filter_firBlock_left_add_225_carry[23]), .YC(my_FIR_filter_firBlock_left_add_225_carry[24]), .YS(my_FIR_filter_firBlock_left_N184));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_24 ( .A(n395),  .B(my_FIR_filter_firBlock_left_multProducts[56]),  .C(my_FIR_filter_firBlock_left_add_225_carry[24]), .YC(my_FIR_filter_firBlock_left_add_225_carry[25]), .YS(my_FIR_filter_firBlock_left_N185));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_25 ( .A(n396),  .B(my_FIR_filter_firBlock_left_multProducts[57]),  .C(my_FIR_filter_firBlock_left_add_225_carry[25]), .YC(my_FIR_filter_firBlock_left_add_225_carry[26]), .YS(my_FIR_filter_firBlock_left_N186));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_26 ( .A(n397),  .B(my_FIR_filter_firBlock_left_multProducts[58]),  .C(my_FIR_filter_firBlock_left_add_225_carry[26]), .YC(my_FIR_filter_firBlock_left_add_225_carry[27]), .YS(my_FIR_filter_firBlock_left_N187));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_27 ( .A(n398),  .B(my_FIR_filter_firBlock_left_multProducts[59]),  .C(my_FIR_filter_firBlock_left_add_225_carry[27]), .YC(my_FIR_filter_firBlock_left_add_225_carry[28]), .YS(my_FIR_filter_firBlock_left_N188));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_28 ( .A(n399),  .B(my_FIR_filter_firBlock_left_multProducts[60]),  .C(my_FIR_filter_firBlock_left_add_225_carry[28]), .YC(my_FIR_filter_firBlock_left_add_225_carry[29]), .YS(my_FIR_filter_firBlock_left_N189));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_29 ( .A(n400),  .B(my_FIR_filter_firBlock_left_multProducts[61]),  .C(my_FIR_filter_firBlock_left_add_225_carry[29]), .YC(my_FIR_filter_firBlock_left_add_225_carry[30]), .YS(my_FIR_filter_firBlock_left_N190));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_30 ( .A(n401),  .B(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[35]),  .C(my_FIR_filter_firBlock_left_add_225_carry[30]), .YC(my_FIR_filter_firBlock_left_add_225_carry[31]), .YS(my_FIR_filter_firBlock_left_N191));
   FAX1 my_FIR_filter_firBlock_left_add_225_U1_31 ( .A(n216),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_225_carry[31]), .YS(my_FIR_filter_firBlock_left_N192));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_1 ( .A(n295),  .B(my_FIR_filter_firBlock_left_multProducts[34]),  .C(n524), .YC(my_FIR_filter_firBlock_left_add_226_carry[2]), .YS(my_FIR_filter_firBlock_left_N194));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_2 ( .A(n187),  .B(my_FIR_filter_firBlock_left_multProducts[35]),  .C(my_FIR_filter_firBlock_left_add_226_carry[2]), .YC(my_FIR_filter_firBlock_left_add_226_carry[3]), .YS(my_FIR_filter_firBlock_left_N195));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_3 ( .A(n188),  .B(my_FIR_filter_firBlock_left_multProducts[36]),  .C(my_FIR_filter_firBlock_left_add_226_carry[3]), .YC(my_FIR_filter_firBlock_left_add_226_carry[4]), .YS(my_FIR_filter_firBlock_left_N196));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_4 ( .A(n189),  .B(my_FIR_filter_firBlock_left_multProducts[37]),  .C(my_FIR_filter_firBlock_left_add_226_carry[4]), .YC(my_FIR_filter_firBlock_left_add_226_carry[5]), .YS(my_FIR_filter_firBlock_left_N197));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_5 ( .A(n190),  .B(my_FIR_filter_firBlock_left_multProducts[38]),  .C(my_FIR_filter_firBlock_left_add_226_carry[5]), .YC(my_FIR_filter_firBlock_left_add_226_carry[6]), .YS(my_FIR_filter_firBlock_left_N198));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_6 ( .A(n191),  .B(my_FIR_filter_firBlock_left_multProducts[39]),  .C(my_FIR_filter_firBlock_left_add_226_carry[6]), .YC(my_FIR_filter_firBlock_left_add_226_carry[7]), .YS(my_FIR_filter_firBlock_left_N199));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_7 ( .A(n192),  .B(my_FIR_filter_firBlock_left_multProducts[40]),  .C(my_FIR_filter_firBlock_left_add_226_carry[7]), .YC(my_FIR_filter_firBlock_left_add_226_carry[8]), .YS(my_FIR_filter_firBlock_left_N200));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_8 ( .A(n193),  .B(my_FIR_filter_firBlock_left_multProducts[41]),  .C(my_FIR_filter_firBlock_left_add_226_carry[8]), .YC(my_FIR_filter_firBlock_left_add_226_carry[9]), .YS(my_FIR_filter_firBlock_left_N201));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_9 ( .A(n194),  .B(my_FIR_filter_firBlock_left_multProducts[42]),  .C(my_FIR_filter_firBlock_left_add_226_carry[9]), .YC(my_FIR_filter_firBlock_left_add_226_carry[10]), .YS(my_FIR_filter_firBlock_left_N202));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_10 ( .A(n195),  .B(my_FIR_filter_firBlock_left_multProducts[43]),  .C(my_FIR_filter_firBlock_left_add_226_carry[10]), .YC(my_FIR_filter_firBlock_left_add_226_carry[11]), .YS(my_FIR_filter_firBlock_left_N203));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_11 ( .A(n196),  .B(my_FIR_filter_firBlock_left_multProducts[44]),  .C(my_FIR_filter_firBlock_left_add_226_carry[11]), .YC(my_FIR_filter_firBlock_left_add_226_carry[12]), .YS(my_FIR_filter_firBlock_left_N204));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_12 ( .A(n197),  .B(my_FIR_filter_firBlock_left_multProducts[45]),  .C(my_FIR_filter_firBlock_left_add_226_carry[12]), .YC(my_FIR_filter_firBlock_left_add_226_carry[13]), .YS(my_FIR_filter_firBlock_left_N205));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_13 ( .A(n198),  .B(my_FIR_filter_firBlock_left_multProducts[46]),  .C(my_FIR_filter_firBlock_left_add_226_carry[13]), .YC(my_FIR_filter_firBlock_left_add_226_carry[14]), .YS(my_FIR_filter_firBlock_left_N206));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_14 ( .A(n199),  .B(my_FIR_filter_firBlock_left_multProducts[47]),  .C(my_FIR_filter_firBlock_left_add_226_carry[14]), .YC(my_FIR_filter_firBlock_left_add_226_carry[15]), .YS(my_FIR_filter_firBlock_left_N207));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_15 ( .A(n200),  .B(my_FIR_filter_firBlock_left_multProducts[48]),  .C(my_FIR_filter_firBlock_left_add_226_carry[15]), .YC(my_FIR_filter_firBlock_left_add_226_carry[16]), .YS(my_FIR_filter_firBlock_left_N208));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_16 ( .A(n201),  .B(my_FIR_filter_firBlock_left_multProducts[49]),  .C(my_FIR_filter_firBlock_left_add_226_carry[16]), .YC(my_FIR_filter_firBlock_left_add_226_carry[17]), .YS(my_FIR_filter_firBlock_left_N209));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_17 ( .A(n202),  .B(my_FIR_filter_firBlock_left_multProducts[50]),  .C(my_FIR_filter_firBlock_left_add_226_carry[17]), .YC(my_FIR_filter_firBlock_left_add_226_carry[18]), .YS(my_FIR_filter_firBlock_left_N210));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_18 ( .A(n203),  .B(my_FIR_filter_firBlock_left_multProducts[51]),  .C(my_FIR_filter_firBlock_left_add_226_carry[18]), .YC(my_FIR_filter_firBlock_left_add_226_carry[19]), .YS(my_FIR_filter_firBlock_left_N211));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_19 ( .A(n204),  .B(my_FIR_filter_firBlock_left_multProducts[52]),  .C(my_FIR_filter_firBlock_left_add_226_carry[19]), .YC(my_FIR_filter_firBlock_left_add_226_carry[20]), .YS(my_FIR_filter_firBlock_left_N212));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_20 ( .A(n205),  .B(my_FIR_filter_firBlock_left_multProducts[53]),  .C(my_FIR_filter_firBlock_left_add_226_carry[20]), .YC(my_FIR_filter_firBlock_left_add_226_carry[21]), .YS(my_FIR_filter_firBlock_left_N213));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_21 ( .A(n206),  .B(my_FIR_filter_firBlock_left_multProducts[54]),  .C(my_FIR_filter_firBlock_left_add_226_carry[21]), .YC(my_FIR_filter_firBlock_left_add_226_carry[22]), .YS(my_FIR_filter_firBlock_left_N214));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_22 ( .A(n207),  .B(my_FIR_filter_firBlock_left_multProducts[55]),  .C(my_FIR_filter_firBlock_left_add_226_carry[22]), .YC(my_FIR_filter_firBlock_left_add_226_carry[23]), .YS(my_FIR_filter_firBlock_left_N215));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_23 ( .A(n208),  .B(my_FIR_filter_firBlock_left_multProducts[56]),  .C(my_FIR_filter_firBlock_left_add_226_carry[23]), .YC(my_FIR_filter_firBlock_left_add_226_carry[24]), .YS(my_FIR_filter_firBlock_left_N216));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_24 ( .A(n209),  .B(my_FIR_filter_firBlock_left_multProducts[57]),  .C(my_FIR_filter_firBlock_left_add_226_carry[24]), .YC(my_FIR_filter_firBlock_left_add_226_carry[25]), .YS(my_FIR_filter_firBlock_left_N217));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_25 ( .A(n210),  .B(my_FIR_filter_firBlock_left_multProducts[58]),  .C(my_FIR_filter_firBlock_left_add_226_carry[25]), .YC(my_FIR_filter_firBlock_left_add_226_carry[26]), .YS(my_FIR_filter_firBlock_left_N218));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_26 ( .A(n211),  .B(my_FIR_filter_firBlock_left_multProducts[59]),  .C(my_FIR_filter_firBlock_left_add_226_carry[26]), .YC(my_FIR_filter_firBlock_left_add_226_carry[27]), .YS(my_FIR_filter_firBlock_left_N219));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_27 ( .A(n212),  .B(my_FIR_filter_firBlock_left_multProducts[60]),  .C(my_FIR_filter_firBlock_left_add_226_carry[27]), .YC(my_FIR_filter_firBlock_left_add_226_carry[28]), .YS(my_FIR_filter_firBlock_left_N220));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_28 ( .A(n213),  .B(my_FIR_filter_firBlock_left_multProducts[61]),  .C(my_FIR_filter_firBlock_left_add_226_carry[28]), .YC(my_FIR_filter_firBlock_left_add_226_carry[29]), .YS(my_FIR_filter_firBlock_left_N221));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_29 ( .A(n214),  .B(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[35]),  .C(my_FIR_filter_firBlock_left_add_226_carry[29]), .YC(my_FIR_filter_firBlock_left_add_226_carry[30]), .YS(my_FIR_filter_firBlock_left_N222));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_30 ( .A(n215),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_226_carry[30]), .YC(my_FIR_filter_firBlock_left_add_226_carry[31]), .YS(my_FIR_filter_firBlock_left_N223));
   FAX1 my_FIR_filter_firBlock_left_add_226_U1_31 ( .A(n119),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_226_carry[31]), .YS(my_FIR_filter_firBlock_left_N224));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_1 ( .A(n464),  .B(my_FIR_filter_firBlock_left_multProducts[63]),  .C(n525), .YC(my_FIR_filter_firBlock_left_add_227_carry[2]), .YS(my_FIR_filter_firBlock_left_N226));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_2 ( .A(n345),  .B(my_FIR_filter_firBlock_left_multProducts[64]),  .C(my_FIR_filter_firBlock_left_add_227_carry[2]), .YC(my_FIR_filter_firBlock_left_add_227_carry[3]), .YS(my_FIR_filter_firBlock_left_N227));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_3 ( .A(n346),  .B(my_FIR_filter_firBlock_left_multProducts[65]),  .C(my_FIR_filter_firBlock_left_add_227_carry[3]), .YC(my_FIR_filter_firBlock_left_add_227_carry[4]), .YS(my_FIR_filter_firBlock_left_N228));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_4 ( .A(n347),  .B(my_FIR_filter_firBlock_left_multProducts[66]),  .C(my_FIR_filter_firBlock_left_add_227_carry[4]), .YC(my_FIR_filter_firBlock_left_add_227_carry[5]), .YS(my_FIR_filter_firBlock_left_N229));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_5 ( .A(n348),  .B(my_FIR_filter_firBlock_left_multProducts[67]),  .C(my_FIR_filter_firBlock_left_add_227_carry[5]), .YC(my_FIR_filter_firBlock_left_add_227_carry[6]), .YS(my_FIR_filter_firBlock_left_N230));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_6 ( .A(n349),  .B(my_FIR_filter_firBlock_left_multProducts[68]),  .C(my_FIR_filter_firBlock_left_add_227_carry[6]), .YC(my_FIR_filter_firBlock_left_add_227_carry[7]), .YS(my_FIR_filter_firBlock_left_N231));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_7 ( .A(n350),  .B(my_FIR_filter_firBlock_left_multProducts[69]),  .C(my_FIR_filter_firBlock_left_add_227_carry[7]), .YC(my_FIR_filter_firBlock_left_add_227_carry[8]), .YS(my_FIR_filter_firBlock_left_N232));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_8 ( .A(n351),  .B(my_FIR_filter_firBlock_left_multProducts[70]),  .C(my_FIR_filter_firBlock_left_add_227_carry[8]), .YC(my_FIR_filter_firBlock_left_add_227_carry[9]), .YS(my_FIR_filter_firBlock_left_N233));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_9 ( .A(n352),  .B(my_FIR_filter_firBlock_left_multProducts[71]),  .C(my_FIR_filter_firBlock_left_add_227_carry[9]), .YC(my_FIR_filter_firBlock_left_add_227_carry[10]), .YS(my_FIR_filter_firBlock_left_N234));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_10 ( .A(n353),  .B(my_FIR_filter_firBlock_left_multProducts[72]),  .C(my_FIR_filter_firBlock_left_add_227_carry[10]), .YC(my_FIR_filter_firBlock_left_add_227_carry[11]), .YS(my_FIR_filter_firBlock_left_N235));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_11 ( .A(n354),  .B(my_FIR_filter_firBlock_left_multProducts[73]),  .C(my_FIR_filter_firBlock_left_add_227_carry[11]), .YC(my_FIR_filter_firBlock_left_add_227_carry[12]), .YS(my_FIR_filter_firBlock_left_N236));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_12 ( .A(n355),  .B(my_FIR_filter_firBlock_left_multProducts[74]),  .C(my_FIR_filter_firBlock_left_add_227_carry[12]), .YC(my_FIR_filter_firBlock_left_add_227_carry[13]), .YS(my_FIR_filter_firBlock_left_N237));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_13 ( .A(n356),  .B(my_FIR_filter_firBlock_left_multProducts[75]),  .C(my_FIR_filter_firBlock_left_add_227_carry[13]), .YC(my_FIR_filter_firBlock_left_add_227_carry[14]), .YS(my_FIR_filter_firBlock_left_N238));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_14 ( .A(n357),  .B(my_FIR_filter_firBlock_left_multProducts[76]),  .C(my_FIR_filter_firBlock_left_add_227_carry[14]), .YC(my_FIR_filter_firBlock_left_add_227_carry[15]), .YS(my_FIR_filter_firBlock_left_N239));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_15 ( .A(n358),  .B(my_FIR_filter_firBlock_left_multProducts[77]),  .C(my_FIR_filter_firBlock_left_add_227_carry[15]), .YC(my_FIR_filter_firBlock_left_add_227_carry[16]), .YS(my_FIR_filter_firBlock_left_N240));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_16 ( .A(n359),  .B(my_FIR_filter_firBlock_left_multProducts[78]),  .C(my_FIR_filter_firBlock_left_add_227_carry[16]), .YC(my_FIR_filter_firBlock_left_add_227_carry[17]), .YS(my_FIR_filter_firBlock_left_N241));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_17 ( .A(n360),  .B(my_FIR_filter_firBlock_left_multProducts[79]),  .C(my_FIR_filter_firBlock_left_add_227_carry[17]), .YC(my_FIR_filter_firBlock_left_add_227_carry[18]), .YS(my_FIR_filter_firBlock_left_N242));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_18 ( .A(n361),  .B(my_FIR_filter_firBlock_left_multProducts[80]),  .C(my_FIR_filter_firBlock_left_add_227_carry[18]), .YC(my_FIR_filter_firBlock_left_add_227_carry[19]), .YS(my_FIR_filter_firBlock_left_N243));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_19 ( .A(n362),  .B(my_FIR_filter_firBlock_left_multProducts[81]),  .C(my_FIR_filter_firBlock_left_add_227_carry[19]), .YC(my_FIR_filter_firBlock_left_add_227_carry[20]), .YS(my_FIR_filter_firBlock_left_N244));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_20 ( .A(n363),  .B(my_FIR_filter_firBlock_left_multProducts[82]),  .C(my_FIR_filter_firBlock_left_add_227_carry[20]), .YC(my_FIR_filter_firBlock_left_add_227_carry[21]), .YS(my_FIR_filter_firBlock_left_N245));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_21 ( .A(n364),  .B(my_FIR_filter_firBlock_left_multProducts[83]),  .C(my_FIR_filter_firBlock_left_add_227_carry[21]), .YC(my_FIR_filter_firBlock_left_add_227_carry[22]), .YS(my_FIR_filter_firBlock_left_N246));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_22 ( .A(n365),  .B(my_FIR_filter_firBlock_left_multProducts[84]),  .C(my_FIR_filter_firBlock_left_add_227_carry[22]), .YC(my_FIR_filter_firBlock_left_add_227_carry[23]), .YS(my_FIR_filter_firBlock_left_N247));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_23 ( .A(n366),  .B(my_FIR_filter_firBlock_left_multProducts[85]),  .C(my_FIR_filter_firBlock_left_add_227_carry[23]), .YC(my_FIR_filter_firBlock_left_add_227_carry[24]), .YS(my_FIR_filter_firBlock_left_N248));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_24 ( .A(n367),  .B(my_FIR_filter_firBlock_left_multProducts[86]),  .C(my_FIR_filter_firBlock_left_add_227_carry[24]), .YC(my_FIR_filter_firBlock_left_add_227_carry[25]), .YS(my_FIR_filter_firBlock_left_N249));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_25 ( .A(n368),  .B(my_FIR_filter_firBlock_left_multProducts[87]),  .C(my_FIR_filter_firBlock_left_add_227_carry[25]), .YC(my_FIR_filter_firBlock_left_add_227_carry[26]), .YS(my_FIR_filter_firBlock_left_N250));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_26 ( .A(n369),  .B(my_FIR_filter_firBlock_left_multProducts[88]),  .C(my_FIR_filter_firBlock_left_add_227_carry[26]), .YC(my_FIR_filter_firBlock_left_add_227_carry[27]), .YS(my_FIR_filter_firBlock_left_N251));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_27 ( .A(n370),  .B(my_FIR_filter_firBlock_left_multProducts[89]),  .C(my_FIR_filter_firBlock_left_add_227_carry[27]), .YC(my_FIR_filter_firBlock_left_add_227_carry[28]), .YS(my_FIR_filter_firBlock_left_N252));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_28 ( .A(n371),  .B(my_FIR_filter_firBlock_left_multProducts[90]),  .C(my_FIR_filter_firBlock_left_add_227_carry[28]), .YC(my_FIR_filter_firBlock_left_add_227_carry[29]), .YS(my_FIR_filter_firBlock_left_N253));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_29 ( .A(n372),  .B(my_FIR_filter_firBlock_left_multProducts[90]),  .C(my_FIR_filter_firBlock_left_add_227_carry[29]), .YC(my_FIR_filter_firBlock_left_add_227_carry[30]), .YS(my_FIR_filter_firBlock_left_N254));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_30 ( .A(n118),  .B(my_FIR_filter_firBlock_left_multProducts[90]),  .C(my_FIR_filter_firBlock_left_add_227_carry[30]), .YC(my_FIR_filter_firBlock_left_add_227_carry[31]), .YS(my_FIR_filter_firBlock_left_N255));
   FAX1 my_FIR_filter_firBlock_left_add_227_U1_31 ( .A(n186),  .B(my_FIR_filter_firBlock_left_multProducts[90]),  .C(my_FIR_filter_firBlock_left_add_227_carry[31]), .YS(my_FIR_filter_firBlock_left_N256));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_1 ( .A(n294),  .B(n485),  .C(n516), .YC(my_FIR_filter_firBlock_left_add_228_carry[2]), .YS(my_FIR_filter_firBlock_left_N258));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_2 ( .A(n169),  .B(n483),  .C(my_FIR_filter_firBlock_left_add_228_carry[2]), .YC(my_FIR_filter_firBlock_left_add_228_carry[3]), .YS(my_FIR_filter_firBlock_left_N259));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_3 ( .A(n170),  .B(n484),  .C(my_FIR_filter_firBlock_left_add_228_carry[3]), .YC(my_FIR_filter_firBlock_left_add_228_carry[4]), .YS(my_FIR_filter_firBlock_left_N260));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_4 ( .A(n171),  .B(n482),  .C(my_FIR_filter_firBlock_left_add_228_carry[4]), .YC(my_FIR_filter_firBlock_left_add_228_carry[5]), .YS(my_FIR_filter_firBlock_left_N261));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_5 ( .A(n105),  .B(n316),  .C(my_FIR_filter_firBlock_left_add_228_carry[5]), .YC(my_FIR_filter_firBlock_left_add_228_carry[6]), .YS(my_FIR_filter_firBlock_left_N262));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_6 ( .A(n106),  .B(n315),  .C(my_FIR_filter_firBlock_left_add_228_carry[6]), .YC(my_FIR_filter_firBlock_left_add_228_carry[7]), .YS(my_FIR_filter_firBlock_left_N263));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_7 ( .A(n107),  .B(n314),  .C(my_FIR_filter_firBlock_left_add_228_carry[7]), .YC(my_FIR_filter_firBlock_left_add_228_carry[8]), .YS(my_FIR_filter_firBlock_left_N264));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_8 ( .A(n108),  .B(n313),  .C(my_FIR_filter_firBlock_left_add_228_carry[8]), .YC(my_FIR_filter_firBlock_left_add_228_carry[9]), .YS(my_FIR_filter_firBlock_left_N265));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_9 ( .A(n172),  .B(n481),  .C(my_FIR_filter_firBlock_left_add_228_carry[9]), .YC(my_FIR_filter_firBlock_left_add_228_carry[10]), .YS(my_FIR_filter_firBlock_left_N266));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_10 ( .A(n173),  .B(n480),  .C(my_FIR_filter_firBlock_left_add_228_carry[10]), .YC(my_FIR_filter_firBlock_left_add_228_carry[11]), .YS(my_FIR_filter_firBlock_left_N267));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_11 ( .A(n174),  .B(n479),  .C(my_FIR_filter_firBlock_left_add_228_carry[11]), .YC(my_FIR_filter_firBlock_left_add_228_carry[12]), .YS(my_FIR_filter_firBlock_left_N268));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_12 ( .A(n175),  .B(n478),  .C(my_FIR_filter_firBlock_left_add_228_carry[12]), .YC(my_FIR_filter_firBlock_left_add_228_carry[13]), .YS(my_FIR_filter_firBlock_left_N269));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_13 ( .A(n109),  .B(n312),  .C(my_FIR_filter_firBlock_left_add_228_carry[13]), .YC(my_FIR_filter_firBlock_left_add_228_carry[14]), .YS(my_FIR_filter_firBlock_left_N270));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_14 ( .A(n110),  .B(n311),  .C(my_FIR_filter_firBlock_left_add_228_carry[14]), .YC(my_FIR_filter_firBlock_left_add_228_carry[15]), .YS(my_FIR_filter_firBlock_left_N271));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_15 ( .A(n111),  .B(n310),  .C(my_FIR_filter_firBlock_left_add_228_carry[15]), .YC(my_FIR_filter_firBlock_left_add_228_carry[16]), .YS(my_FIR_filter_firBlock_left_N272));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_16 ( .A(n112),  .B(n309),  .C(my_FIR_filter_firBlock_left_add_228_carry[16]), .YC(my_FIR_filter_firBlock_left_add_228_carry[17]), .YS(my_FIR_filter_firBlock_left_N273));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_17 ( .A(n176),  .B(n477),  .C(my_FIR_filter_firBlock_left_add_228_carry[17]), .YC(my_FIR_filter_firBlock_left_add_228_carry[18]), .YS(my_FIR_filter_firBlock_left_N274));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_18 ( .A(n177),  .B(n476),  .C(my_FIR_filter_firBlock_left_add_228_carry[18]), .YC(my_FIR_filter_firBlock_left_add_228_carry[19]), .YS(my_FIR_filter_firBlock_left_N275));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_19 ( .A(n178),  .B(n475),  .C(my_FIR_filter_firBlock_left_add_228_carry[19]), .YC(my_FIR_filter_firBlock_left_add_228_carry[20]), .YS(my_FIR_filter_firBlock_left_N276));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_20 ( .A(n179),  .B(n474),  .C(my_FIR_filter_firBlock_left_add_228_carry[20]), .YC(my_FIR_filter_firBlock_left_add_228_carry[21]), .YS(my_FIR_filter_firBlock_left_N277));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_21 ( .A(n113),  .B(n308),  .C(my_FIR_filter_firBlock_left_add_228_carry[21]), .YC(my_FIR_filter_firBlock_left_add_228_carry[22]), .YS(my_FIR_filter_firBlock_left_N278));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_22 ( .A(n114),  .B(n307),  .C(my_FIR_filter_firBlock_left_add_228_carry[22]), .YC(my_FIR_filter_firBlock_left_add_228_carry[23]), .YS(my_FIR_filter_firBlock_left_N279));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_23 ( .A(n115),  .B(n306),  .C(my_FIR_filter_firBlock_left_add_228_carry[23]), .YC(my_FIR_filter_firBlock_left_add_228_carry[24]), .YS(my_FIR_filter_firBlock_left_N280));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_24 ( .A(n116),  .B(n305),  .C(my_FIR_filter_firBlock_left_add_228_carry[24]), .YC(my_FIR_filter_firBlock_left_add_228_carry[25]), .YS(my_FIR_filter_firBlock_left_N281));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_25 ( .A(n180),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_228_carry[25]), .YC(my_FIR_filter_firBlock_left_add_228_carry[26]), .YS(my_FIR_filter_firBlock_left_N282));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_26 ( .A(n181),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_228_carry[26]), .YC(my_FIR_filter_firBlock_left_add_228_carry[27]), .YS(my_FIR_filter_firBlock_left_N283));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_27 ( .A(n182),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_228_carry[27]), .YC(my_FIR_filter_firBlock_left_add_228_carry[28]), .YS(my_FIR_filter_firBlock_left_N284));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_28 ( .A(n183),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_228_carry[28]), .YC(my_FIR_filter_firBlock_left_add_228_carry[29]), .YS(my_FIR_filter_firBlock_left_N285));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_29 ( .A(n184),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_228_carry[29]), .YC(my_FIR_filter_firBlock_left_add_228_carry[30]), .YS(my_FIR_filter_firBlock_left_N286));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_30 ( .A(n185),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_228_carry[30]), .YC(my_FIR_filter_firBlock_left_add_228_carry[31]), .YS(my_FIR_filter_firBlock_left_N287));
   FAX1 my_FIR_filter_firBlock_left_add_228_U1_31 ( .A(n117),  .B(n486),  .C(my_FIR_filter_firBlock_left_add_228_carry[31]), .YS(my_FIR_filter_firBlock_left_N288));
   FAX1 add_63_U1_1 ( .A(n463),  .B(n104),  .C(n526), .YC(add_63_carry[2]), .YS(outData_in[1]));
   FAX1 add_63_U1_2 ( .A(n344),  .B(n139),  .C(add_63_carry[2]), .YC(add_63_carry[3]), .YS(outData_in[2]));
   FAX1 add_63_U1_3 ( .A(n343),  .B(n140),  .C(add_63_carry[3]), .YC(add_63_carry[4]), .YS(outData_in[3]));
   FAX1 add_63_U1_4 ( .A(n342),  .B(n141),  .C(add_63_carry[4]), .YC(add_63_carry[5]), .YS(outData_in[4]));
   FAX1 add_63_U1_5 ( .A(n341),  .B(n142),  .C(add_63_carry[5]), .YC(add_63_carry[6]), .YS(outData_in[5]));
   FAX1 add_63_U1_6 ( .A(n340),  .B(n143),  .C(add_63_carry[6]), .YC(add_63_carry[7]), .YS(outData_in[6]));
   FAX1 add_63_U1_7 ( .A(n339),  .B(n144),  .C(add_63_carry[7]), .YC(add_63_carry[8]), .YS(outData_in[7]));
   FAX1 add_63_U1_8 ( .A(n338),  .B(n145),  .C(add_63_carry[8]), .YC(add_63_carry[9]), .YS(outData_in[8]));
   FAX1 add_63_U1_9 ( .A(n337),  .B(n146),  .C(add_63_carry[9]), .YC(add_63_carry[10]), .YS(outData_in[9]));
   FAX1 add_63_U1_10 ( .A(n336),  .B(n147),  .C(add_63_carry[10]), .YC(add_63_carry[11]), .YS(outData_in[10]));
   FAX1 add_63_U1_11 ( .A(n335),  .B(n148),  .C(add_63_carry[11]), .YC(add_63_carry[12]), .YS(outData_in[11]));
   FAX1 add_63_U1_12 ( .A(n334),  .B(n149),  .C(add_63_carry[12]), .YC(add_63_carry[13]), .YS(outData_in[12]));
   FAX1 add_63_U1_13 ( .A(n333),  .B(n150),  .C(add_63_carry[13]), .YC(add_63_carry[14]), .YS(outData_in[13]));
   FAX1 add_63_U1_14 ( .A(n332),  .B(n151),  .C(add_63_carry[14]), .YC(add_63_carry[15]), .YS(outData_in[14]));
   FAX1 add_63_U1_15 ( .A(n331),  .B(n152),  .C(add_63_carry[15]), .YC(add_63_carry[16]), .YS(outData_in[15]));
   FAX1 add_63_U1_16 ( .A(n330),  .B(n153),  .C(add_63_carry[16]), .YC(add_63_carry[17]), .YS(outData_in[16]));
   FAX1 add_63_U1_17 ( .A(n329),  .B(n154),  .C(add_63_carry[17]), .YC(add_63_carry[18]), .YS(outData_in[17]));
   FAX1 add_63_U1_18 ( .A(n328),  .B(n155),  .C(add_63_carry[18]), .YC(add_63_carry[19]), .YS(outData_in[18]));
   FAX1 add_63_U1_19 ( .A(n327),  .B(n156),  .C(add_63_carry[19]), .YC(add_63_carry[20]), .YS(outData_in[19]));
   FAX1 add_63_U1_20 ( .A(n326),  .B(n157),  .C(add_63_carry[20]), .YC(add_63_carry[21]), .YS(outData_in[20]));
   FAX1 add_63_U1_21 ( .A(n325),  .B(n158),  .C(add_63_carry[21]), .YC(add_63_carry[22]), .YS(outData_in[21]));
   FAX1 add_63_U1_22 ( .A(n324),  .B(n159),  .C(add_63_carry[22]), .YC(add_63_carry[23]), .YS(outData_in[22]));
   FAX1 add_63_U1_23 ( .A(n323),  .B(n160),  .C(add_63_carry[23]), .YC(add_63_carry[24]), .YS(outData_in[23]));
   FAX1 add_63_U1_24 ( .A(n322),  .B(n161),  .C(add_63_carry[24]), .YC(add_63_carry[25]), .YS(outData_in[24]));
   FAX1 add_63_U1_25 ( .A(n321),  .B(n162),  .C(add_63_carry[25]), .YC(add_63_carry[26]), .YS(outData_in[25]));
   FAX1 add_63_U1_26 ( .A(n320),  .B(n163),  .C(add_63_carry[26]), .YC(add_63_carry[27]), .YS(outData_in[26]));
   FAX1 add_63_U1_27 ( .A(n460),  .B(n166),  .C(add_63_carry[27]), .YC(add_63_carry[28]), .YS(outData_in[27]));
   FAX1 add_63_U1_28 ( .A(n462),  .B(n167),  .C(add_63_carry[28]), .YC(add_63_carry[29]), .YS(outData_in[28]));
   FAX1 add_63_U1_29 ( .A(n461),  .B(n168),  .C(add_63_carry[29]), .YC(add_63_carry[30]), .YS(outData_in[29]));
   FAX1 add_63_U1_30 ( .A(n319),  .B(n164),  .C(add_63_carry[30]), .YC(add_63_carry[31]), .YS(outData_in[30]));
   FAX1 add_63_U1_31 ( .A(n318),  .B(n165),  .C(add_63_carry[31]), .YS(outData_in[31]));
   AND2X1 U68 ( .A(n103),  .B(n138), .Y(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[5]));
   AND2X1 U69 ( .A(my_FIR_filter_firBlock_left_multProducts[62]),  .B(n136), .Y(n518));
   AND2X1 U70 ( .A(my_FIR_filter_firBlock_left_multProducts[33]),  .B(n472), .Y(n519));
   AND2X1 U71 ( .A(my_FIR_filter_firBlock_left_multProducts[32]),  .B(n302), .Y(n520));
   AND2X1 U72 ( .A(my_FIR_filter_firBlock_left_multProducts[0]),  .B(n471), .Y(n521));
   AND2X1 U73 ( .A(my_FIR_filter_firBlock_left_multProducts[0]),  .B(n301), .Y(n522));
   AND2X1 U74 ( .A(my_FIR_filter_firBlock_left_multProducts[32]),  .B(n470), .Y(n523));
   AND2X1 U75 ( .A(my_FIR_filter_firBlock_left_multProducts[33]),  .B(n300), .Y(n524));
   AND2X1 U76 ( .A(my_FIR_filter_firBlock_left_multProducts[62]),  .B(n469), .Y(n525));
   AND2X1 U77 ( .A(n317),  .B(n135), .Y(n516));
   AND2X1 U78 ( .A(n468),  .B(n299), .Y(n526));
   XNOR2X1 U79 ( .A(n572),  .B(n573), .Y(n66));
   BUFX2 U80 ( .A(my_FIR_filter_firBlock_left_firStep[30]), .Y(puf_52_wire_1));
   BUFX2 U81 ( .A(my_FIR_filter_firBlock_left_firStep[29]), .Y(puf_53_wire_1));
   BUFX2 U82 ( .A(my_FIR_filter_firBlock_left_firStep[28]), .Y(puf_54_wire_1));
   BUFX2 U83 ( .A(my_FIR_filter_firBlock_left_firStep[27]), .Y(puf_55_wire_1));
   BUFX2 U84 ( .A(my_FIR_filter_firBlock_left_firStep[26]), .Y(puf_56_wire_1));
   BUFX2 U85 ( .A(my_FIR_filter_firBlock_left_firStep[25]), .Y(puf_57_wire_1));
   BUFX2 U86 ( .A(my_FIR_filter_firBlock_left_firStep[24]), .Y(puf_58_wire_1));
   BUFX2 U87 ( .A(my_FIR_filter_firBlock_left_firStep[23]), .Y(puf_59_wire_1));
   BUFX2 U88 ( .A(my_FIR_filter_firBlock_left_firStep[22]), .Y(puf_60_wire_1));
   BUFX2 U89 ( .A(my_FIR_filter_firBlock_left_firStep[21]), .Y(puf_61_wire_1));
   BUFX2 U90 ( .A(my_FIR_filter_firBlock_left_firStep[20]), .Y(puf_62_wire_1));
   BUFX2 U91 ( .A(my_FIR_filter_firBlock_left_firStep[19]), .Y(puf_63_wire_1));
   BUFX2 U92 ( .A(my_FIR_filter_firBlock_left_firStep[18]), .Y(puf_64_wire_1));
   BUFX2 U93 ( .A(my_FIR_filter_firBlock_left_firStep[17]), .Y(puf_65_wire_1));
   BUFX2 U94 ( .A(my_FIR_filter_firBlock_left_firStep[16]), .Y(puf_66_wire_1));
   BUFX2 U95 ( .A(my_FIR_filter_firBlock_left_firStep[15]), .Y(puf_67_wire_1));
   BUFX2 U96 ( .A(my_FIR_filter_firBlock_left_firStep[14]), .Y(puf_68_wire_1));
   BUFX2 U97 ( .A(my_FIR_filter_firBlock_left_firStep[13]), .Y(puf_69_wire_1));
   BUFX2 U98 ( .A(my_FIR_filter_firBlock_left_firStep[12]), .Y(puf_70_wire_1));
   BUFX2 U99 ( .A(my_FIR_filter_firBlock_left_firStep[11]), .Y(puf_71_wire_1));
   BUFX2 U100 ( .A(my_FIR_filter_firBlock_left_firStep[10]), .Y(puf_72_wire_1));
   BUFX2 U101 ( .A(my_FIR_filter_firBlock_left_firStep[9]), .Y(puf_73_wire_1));
   BUFX2 U102 ( .A(my_FIR_filter_firBlock_left_firStep[8]), .Y(puf_74_wire_1));
   BUFX2 U103 ( .A(my_FIR_filter_firBlock_left_firStep[7]), .Y(puf_75_wire_1));
   BUFX2 U104 ( .A(my_FIR_filter_firBlock_left_firStep[6]), .Y(puf_76_wire_1));
   BUFX2 U105 ( .A(my_FIR_filter_firBlock_left_firStep[5]), .Y(puf_77_wire_1));
   BUFX2 U106 ( .A(my_FIR_filter_firBlock_left_firStep[4]), .Y(puf_78_wire_1));
   BUFX2 U107 ( .A(my_FIR_filter_firBlock_left_firStep[3]), .Y(puf_79_wire_1));
   BUFX2 U108 ( .A(my_FIR_filter_firBlock_left_firStep[2]), .Y(puf_80_wire_1));
   BUFX2 U109 ( .A(my_FIR_filter_firBlock_left_firStep[1]), .Y(puf_81_wire_1));
   BUFX2 U110 ( .A(my_FIR_filter_firBlock_left_firStep[0]), .Y(puf_82_wire_1));
   BUFX2 U111 ( .A(my_FIR_filter_firBlock_left_Y_in_0_), .Y(puf_83_wire_1));
   BUFX2 U112 ( .A(n530), .Y(n99));
   BUFX2 U113 ( .A(n531), .Y(n100));
   BUFX2 U114 ( .A(n539), .Y(n101));
   AND2X1 U115 ( .A(n538),  .B(n572), .Y(n540));
   INVX1 U116 ( .A(n540), .Y(n102));
   BUFX2 U117 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_6_), .Y(n103));
   AND2X1 U118 ( .A(n575),  .B(n514), .Y(n527));
   BUFX2 U119 ( .A(rightOut[1]), .Y(n104));
   BUFX2 U120 ( .A(my_FIR_filter_firBlock_left_firStep[36]), .Y(n105));
   BUFX2 U121 ( .A(my_FIR_filter_firBlock_left_firStep[37]), .Y(n106));
   BUFX2 U122 ( .A(my_FIR_filter_firBlock_left_firStep[38]), .Y(n107));
   BUFX2 U123 ( .A(my_FIR_filter_firBlock_left_firStep[39]), .Y(n108));
   BUFX2 U124 ( .A(my_FIR_filter_firBlock_left_firStep[44]), .Y(n109));
   BUFX2 U125 ( .A(my_FIR_filter_firBlock_left_firStep[45]), .Y(n110));
   BUFX2 U126 ( .A(my_FIR_filter_firBlock_left_firStep[46]), .Y(n111));
   BUFX2 U127 ( .A(my_FIR_filter_firBlock_left_firStep[47]), .Y(n112));
   BUFX2 U128 ( .A(my_FIR_filter_firBlock_left_firStep[52]), .Y(n113));
   BUFX2 U129 ( .A(my_FIR_filter_firBlock_left_firStep[53]), .Y(n114));
   BUFX2 U130 ( .A(my_FIR_filter_firBlock_left_firStep[54]), .Y(n115));
   BUFX2 U131 ( .A(my_FIR_filter_firBlock_left_firStep[55]), .Y(n116));
   BUFX2 U132 ( .A(my_FIR_filter_firBlock_left_firStep[62]), .Y(n117));
   BUFX2 U133 ( .A(my_FIR_filter_firBlock_left_firStep[93]), .Y(n118));
   BUFX2 U134 ( .A(my_FIR_filter_firBlock_left_firStep[126]), .Y(n119));
   BUFX2 U135 ( .A(my_FIR_filter_firBlock_left_firStep[222]), .Y(n120));
   BUFX2 U136 ( .A(my_FIR_filter_firBlock_left_firStep[285]), .Y(n121));
   BUFX2 U137 ( .A(my_FIR_filter_firBlock_left_firStep[286]), .Y(n122));
   BUFX2 U138 ( .A(my_FIR_filter_firBlock_left_firStep[292]), .Y(n123));
   BUFX2 U139 ( .A(my_FIR_filter_firBlock_left_firStep[293]), .Y(n124));
   BUFX2 U140 ( .A(my_FIR_filter_firBlock_left_firStep[294]), .Y(n125));
   BUFX2 U141 ( .A(my_FIR_filter_firBlock_left_firStep[295]), .Y(n126));
   BUFX2 U142 ( .A(my_FIR_filter_firBlock_left_firStep[300]), .Y(n127));
   BUFX2 U143 ( .A(my_FIR_filter_firBlock_left_firStep[301]), .Y(n128));
   BUFX2 U144 ( .A(my_FIR_filter_firBlock_left_firStep[302]), .Y(n129));
   BUFX2 U145 ( .A(my_FIR_filter_firBlock_left_firStep[303]), .Y(n130));
   BUFX2 U146 ( .A(my_FIR_filter_firBlock_left_firStep[308]), .Y(n131));
   BUFX2 U147 ( .A(my_FIR_filter_firBlock_left_firStep[309]), .Y(n132));
   BUFX2 U148 ( .A(my_FIR_filter_firBlock_left_firStep[310]), .Y(n133));
   BUFX2 U149 ( .A(my_FIR_filter_firBlock_left_firStep[311]), .Y(n134));
   BUFX2 U150 ( .A(my_FIR_filter_firBlock_left_firStep[31]), .Y(n135));
   BUFX2 U151 ( .A(my_FIR_filter_firBlock_left_firStep[287]), .Y(n136));
   BUFX2 U152 ( .A(inData_in[1]), .Y(n137));
   BUFX2 U153 ( .A(inData_in[4]), .Y(n138));
   BUFX2 U154 ( .A(rightOut[2]), .Y(n139));
   BUFX2 U155 ( .A(rightOut[3]), .Y(n140));
   BUFX2 U156 ( .A(rightOut[4]), .Y(n141));
   BUFX2 U157 ( .A(rightOut[5]), .Y(n142));
   BUFX2 U158 ( .A(rightOut[6]), .Y(n143));
   BUFX2 U159 ( .A(rightOut[7]), .Y(n144));
   BUFX2 U160 ( .A(rightOut[8]), .Y(n145));
   BUFX2 U161 ( .A(rightOut[9]), .Y(n146));
   BUFX2 U162 ( .A(rightOut[10]), .Y(n147));
   BUFX2 U163 ( .A(rightOut[11]), .Y(n148));
   BUFX2 U164 ( .A(rightOut[12]), .Y(n149));
   BUFX2 U165 ( .A(rightOut[13]), .Y(n150));
   BUFX2 U166 ( .A(rightOut[14]), .Y(n151));
   BUFX2 U167 ( .A(rightOut[15]), .Y(n152));
   BUFX2 U168 ( .A(rightOut[16]), .Y(n153));
   BUFX2 U169 ( .A(rightOut[17]), .Y(n154));
   BUFX2 U170 ( .A(rightOut[18]), .Y(n155));
   BUFX2 U171 ( .A(rightOut[19]), .Y(n156));
   BUFX2 U172 ( .A(rightOut[20]), .Y(n157));
   BUFX2 U173 ( .A(rightOut[21]), .Y(n158));
   BUFX2 U174 ( .A(rightOut[22]), .Y(n159));
   BUFX2 U175 ( .A(rightOut[23]), .Y(n160));
   BUFX2 U176 ( .A(rightOut[24]), .Y(n161));
   BUFX2 U177 ( .A(rightOut[25]), .Y(n162));
   BUFX2 U178 ( .A(rightOut[26]), .Y(n163));
   BUFX2 U179 ( .A(rightOut[30]), .Y(n164));
   BUFX2 U180 ( .A(rightOut[31]), .Y(n165));
   BUFX2 U181 ( .A(rightOut[27]), .Y(n166));
   BUFX2 U182 ( .A(rightOut[28]), .Y(n167));
   BUFX2 U183 ( .A(rightOut[29]), .Y(n168));
   BUFX2 U184 ( .A(my_FIR_filter_firBlock_left_firStep[33]), .Y(n169));
   BUFX2 U185 ( .A(my_FIR_filter_firBlock_left_firStep[34]), .Y(n170));
   BUFX2 U186 ( .A(my_FIR_filter_firBlock_left_firStep[35]), .Y(n171));
   BUFX2 U187 ( .A(my_FIR_filter_firBlock_left_firStep[40]), .Y(n172));
   BUFX2 U188 ( .A(my_FIR_filter_firBlock_left_firStep[41]), .Y(n173));
   BUFX2 U189 ( .A(my_FIR_filter_firBlock_left_firStep[42]), .Y(n174));
   BUFX2 U190 ( .A(my_FIR_filter_firBlock_left_firStep[43]), .Y(n175));
   BUFX2 U191 ( .A(my_FIR_filter_firBlock_left_firStep[48]), .Y(n176));
   BUFX2 U192 ( .A(my_FIR_filter_firBlock_left_firStep[49]), .Y(n177));
   BUFX2 U193 ( .A(my_FIR_filter_firBlock_left_firStep[50]), .Y(n178));
   BUFX2 U194 ( .A(my_FIR_filter_firBlock_left_firStep[51]), .Y(n179));
   BUFX2 U195 ( .A(my_FIR_filter_firBlock_left_firStep[56]), .Y(n180));
   BUFX2 U196 ( .A(my_FIR_filter_firBlock_left_firStep[57]), .Y(n181));
   BUFX2 U197 ( .A(my_FIR_filter_firBlock_left_firStep[58]), .Y(n182));
   BUFX2 U198 ( .A(my_FIR_filter_firBlock_left_firStep[59]), .Y(n183));
   BUFX2 U199 ( .A(my_FIR_filter_firBlock_left_firStep[60]), .Y(n184));
   BUFX2 U200 ( .A(my_FIR_filter_firBlock_left_firStep[61]), .Y(n185));
   BUFX2 U201 ( .A(my_FIR_filter_firBlock_left_firStep[94]), .Y(n186));
   BUFX2 U202 ( .A(my_FIR_filter_firBlock_left_firStep[97]), .Y(n187));
   BUFX2 U203 ( .A(my_FIR_filter_firBlock_left_firStep[98]), .Y(n188));
   BUFX2 U204 ( .A(my_FIR_filter_firBlock_left_firStep[99]), .Y(n189));
   BUFX2 U205 ( .A(my_FIR_filter_firBlock_left_firStep[100]), .Y(n190));
   BUFX2 U206 ( .A(my_FIR_filter_firBlock_left_firStep[101]), .Y(n191));
   BUFX2 U207 ( .A(my_FIR_filter_firBlock_left_firStep[102]), .Y(n192));
   BUFX2 U208 ( .A(my_FIR_filter_firBlock_left_firStep[103]), .Y(n193));
   BUFX2 U209 ( .A(my_FIR_filter_firBlock_left_firStep[104]), .Y(n194));
   BUFX2 U210 ( .A(my_FIR_filter_firBlock_left_firStep[105]), .Y(n195));
   BUFX2 U211 ( .A(my_FIR_filter_firBlock_left_firStep[106]), .Y(n196));
   BUFX2 U212 ( .A(my_FIR_filter_firBlock_left_firStep[107]), .Y(n197));
   BUFX2 U213 ( .A(my_FIR_filter_firBlock_left_firStep[108]), .Y(n198));
   BUFX2 U214 ( .A(my_FIR_filter_firBlock_left_firStep[109]), .Y(n199));
   BUFX2 U215 ( .A(my_FIR_filter_firBlock_left_firStep[110]), .Y(n200));
   BUFX2 U216 ( .A(my_FIR_filter_firBlock_left_firStep[111]), .Y(n201));
   BUFX2 U217 ( .A(my_FIR_filter_firBlock_left_firStep[112]), .Y(n202));
   BUFX2 U218 ( .A(my_FIR_filter_firBlock_left_firStep[113]), .Y(n203));
   BUFX2 U219 ( .A(my_FIR_filter_firBlock_left_firStep[114]), .Y(n204));
   BUFX2 U220 ( .A(my_FIR_filter_firBlock_left_firStep[115]), .Y(n205));
   BUFX2 U221 ( .A(my_FIR_filter_firBlock_left_firStep[116]), .Y(n206));
   BUFX2 U222 ( .A(my_FIR_filter_firBlock_left_firStep[117]), .Y(n207));
   BUFX2 U223 ( .A(my_FIR_filter_firBlock_left_firStep[118]), .Y(n208));
   BUFX2 U224 ( .A(my_FIR_filter_firBlock_left_firStep[119]), .Y(n209));
   BUFX2 U225 ( .A(my_FIR_filter_firBlock_left_firStep[120]), .Y(n210));
   BUFX2 U226 ( .A(my_FIR_filter_firBlock_left_firStep[121]), .Y(n211));
   BUFX2 U227 ( .A(my_FIR_filter_firBlock_left_firStep[122]), .Y(n212));
   BUFX2 U228 ( .A(my_FIR_filter_firBlock_left_firStep[123]), .Y(n213));
   BUFX2 U229 ( .A(my_FIR_filter_firBlock_left_firStep[124]), .Y(n214));
   BUFX2 U230 ( .A(my_FIR_filter_firBlock_left_firStep[125]), .Y(n215));
   BUFX2 U231 ( .A(my_FIR_filter_firBlock_left_firStep[158]), .Y(n216));
   BUFX2 U232 ( .A(my_FIR_filter_firBlock_left_firStep[161]), .Y(n217));
   BUFX2 U233 ( .A(my_FIR_filter_firBlock_left_firStep[162]), .Y(n218));
   BUFX2 U234 ( .A(my_FIR_filter_firBlock_left_firStep[163]), .Y(n219));
   BUFX2 U235 ( .A(my_FIR_filter_firBlock_left_firStep[164]), .Y(n220));
   BUFX2 U236 ( .A(my_FIR_filter_firBlock_left_firStep[165]), .Y(n221));
   BUFX2 U237 ( .A(my_FIR_filter_firBlock_left_firStep[166]), .Y(n222));
   BUFX2 U238 ( .A(my_FIR_filter_firBlock_left_firStep[167]), .Y(n223));
   BUFX2 U239 ( .A(my_FIR_filter_firBlock_left_firStep[168]), .Y(n224));
   BUFX2 U240 ( .A(my_FIR_filter_firBlock_left_firStep[169]), .Y(n225));
   BUFX2 U241 ( .A(my_FIR_filter_firBlock_left_firStep[170]), .Y(n226));
   BUFX2 U242 ( .A(my_FIR_filter_firBlock_left_firStep[171]), .Y(n227));
   BUFX2 U243 ( .A(my_FIR_filter_firBlock_left_firStep[172]), .Y(n228));
   BUFX2 U244 ( .A(my_FIR_filter_firBlock_left_firStep[173]), .Y(n229));
   BUFX2 U245 ( .A(my_FIR_filter_firBlock_left_firStep[174]), .Y(n230));
   BUFX2 U246 ( .A(my_FIR_filter_firBlock_left_firStep[175]), .Y(n231));
   BUFX2 U247 ( .A(my_FIR_filter_firBlock_left_firStep[176]), .Y(n232));
   BUFX2 U248 ( .A(my_FIR_filter_firBlock_left_firStep[177]), .Y(n233));
   BUFX2 U249 ( .A(my_FIR_filter_firBlock_left_firStep[178]), .Y(n234));
   BUFX2 U250 ( .A(my_FIR_filter_firBlock_left_firStep[179]), .Y(n235));
   BUFX2 U251 ( .A(my_FIR_filter_firBlock_left_firStep[180]), .Y(n236));
   BUFX2 U252 ( .A(my_FIR_filter_firBlock_left_firStep[181]), .Y(n237));
   BUFX2 U253 ( .A(my_FIR_filter_firBlock_left_firStep[182]), .Y(n238));
   BUFX2 U254 ( .A(my_FIR_filter_firBlock_left_firStep[183]), .Y(n239));
   BUFX2 U255 ( .A(my_FIR_filter_firBlock_left_firStep[184]), .Y(n240));
   BUFX2 U256 ( .A(my_FIR_filter_firBlock_left_firStep[185]), .Y(n241));
   BUFX2 U257 ( .A(my_FIR_filter_firBlock_left_firStep[186]), .Y(n242));
   BUFX2 U258 ( .A(my_FIR_filter_firBlock_left_firStep[187]), .Y(n243));
   BUFX2 U259 ( .A(my_FIR_filter_firBlock_left_firStep[188]), .Y(n244));
   BUFX2 U260 ( .A(my_FIR_filter_firBlock_left_firStep[189]), .Y(n245));
   BUFX2 U261 ( .A(my_FIR_filter_firBlock_left_firStep[225]), .Y(n246));
   BUFX2 U262 ( .A(my_FIR_filter_firBlock_left_firStep[226]), .Y(n247));
   BUFX2 U263 ( .A(my_FIR_filter_firBlock_left_firStep[227]), .Y(n248));
   BUFX2 U264 ( .A(my_FIR_filter_firBlock_left_firStep[228]), .Y(n249));
   BUFX2 U265 ( .A(my_FIR_filter_firBlock_left_firStep[229]), .Y(n250));
   BUFX2 U266 ( .A(my_FIR_filter_firBlock_left_firStep[230]), .Y(n251));
   BUFX2 U267 ( .A(my_FIR_filter_firBlock_left_firStep[231]), .Y(n252));
   BUFX2 U268 ( .A(my_FIR_filter_firBlock_left_firStep[232]), .Y(n253));
   BUFX2 U269 ( .A(my_FIR_filter_firBlock_left_firStep[233]), .Y(n254));
   BUFX2 U270 ( .A(my_FIR_filter_firBlock_left_firStep[234]), .Y(n255));
   BUFX2 U271 ( .A(my_FIR_filter_firBlock_left_firStep[235]), .Y(n256));
   BUFX2 U272 ( .A(my_FIR_filter_firBlock_left_firStep[236]), .Y(n257));
   BUFX2 U273 ( .A(my_FIR_filter_firBlock_left_firStep[237]), .Y(n258));
   BUFX2 U274 ( .A(my_FIR_filter_firBlock_left_firStep[238]), .Y(n259));
   BUFX2 U275 ( .A(my_FIR_filter_firBlock_left_firStep[239]), .Y(n260));
   BUFX2 U276 ( .A(my_FIR_filter_firBlock_left_firStep[240]), .Y(n261));
   BUFX2 U277 ( .A(my_FIR_filter_firBlock_left_firStep[241]), .Y(n262));
   BUFX2 U278 ( .A(my_FIR_filter_firBlock_left_firStep[242]), .Y(n263));
   BUFX2 U279 ( .A(my_FIR_filter_firBlock_left_firStep[243]), .Y(n264));
   BUFX2 U280 ( .A(my_FIR_filter_firBlock_left_firStep[244]), .Y(n265));
   BUFX2 U281 ( .A(my_FIR_filter_firBlock_left_firStep[245]), .Y(n266));
   BUFX2 U282 ( .A(my_FIR_filter_firBlock_left_firStep[246]), .Y(n267));
   BUFX2 U283 ( .A(my_FIR_filter_firBlock_left_firStep[247]), .Y(n268));
   BUFX2 U284 ( .A(my_FIR_filter_firBlock_left_firStep[248]), .Y(n269));
   BUFX2 U285 ( .A(my_FIR_filter_firBlock_left_firStep[249]), .Y(n270));
   BUFX2 U286 ( .A(my_FIR_filter_firBlock_left_firStep[250]), .Y(n271));
   BUFX2 U287 ( .A(my_FIR_filter_firBlock_left_firStep[251]), .Y(n272));
   BUFX2 U288 ( .A(my_FIR_filter_firBlock_left_firStep[252]), .Y(n273));
   BUFX2 U289 ( .A(my_FIR_filter_firBlock_left_firStep[253]), .Y(n274));
   BUFX2 U290 ( .A(my_FIR_filter_firBlock_left_firStep[254]), .Y(n275));
   BUFX2 U291 ( .A(my_FIR_filter_firBlock_left_firStep[289]), .Y(n276));
   BUFX2 U292 ( .A(my_FIR_filter_firBlock_left_firStep[290]), .Y(n277));
   BUFX2 U293 ( .A(my_FIR_filter_firBlock_left_firStep[291]), .Y(n278));
   BUFX2 U294 ( .A(my_FIR_filter_firBlock_left_firStep[296]), .Y(n279));
   BUFX2 U295 ( .A(my_FIR_filter_firBlock_left_firStep[297]), .Y(n280));
   BUFX2 U296 ( .A(my_FIR_filter_firBlock_left_firStep[298]), .Y(n281));
   BUFX2 U297 ( .A(my_FIR_filter_firBlock_left_firStep[299]), .Y(n282));
   BUFX2 U298 ( .A(my_FIR_filter_firBlock_left_firStep[304]), .Y(n283));
   BUFX2 U299 ( .A(my_FIR_filter_firBlock_left_firStep[305]), .Y(n284));
   BUFX2 U300 ( .A(my_FIR_filter_firBlock_left_firStep[306]), .Y(n285));
   BUFX2 U301 ( .A(my_FIR_filter_firBlock_left_firStep[307]), .Y(n286));
   BUFX2 U302 ( .A(my_FIR_filter_firBlock_left_firStep[312]), .Y(n287));
   BUFX2 U303 ( .A(my_FIR_filter_firBlock_left_firStep[313]), .Y(n288));
   BUFX2 U304 ( .A(my_FIR_filter_firBlock_left_firStep[314]), .Y(n289));
   BUFX2 U305 ( .A(my_FIR_filter_firBlock_left_firStep[315]), .Y(n290));
   BUFX2 U306 ( .A(my_FIR_filter_firBlock_left_firStep[316]), .Y(n291));
   BUFX2 U307 ( .A(my_FIR_filter_firBlock_left_firStep[317]), .Y(n292));
   BUFX2 U308 ( .A(my_FIR_filter_firBlock_left_firStep[318]), .Y(n293));
   BUFX2 U309 ( .A(my_FIR_filter_firBlock_left_firStep[32]), .Y(n294));
   BUFX2 U310 ( .A(my_FIR_filter_firBlock_left_firStep[96]), .Y(n295));
   BUFX2 U311 ( .A(my_FIR_filter_firBlock_left_firStep[160]), .Y(n296));
   BUFX2 U312 ( .A(my_FIR_filter_firBlock_left_firStep[224]), .Y(n297));
   BUFX2 U313 ( .A(my_FIR_filter_firBlock_left_firStep[288]), .Y(n298));
   BUFX2 U314 ( .A(rightOut[0]), .Y(n299));
   BUFX2 U315 ( .A(my_FIR_filter_firBlock_left_firStep[95]), .Y(n300));
   BUFX2 U316 ( .A(my_FIR_filter_firBlock_left_firStep[159]), .Y(n301));
   BUFX2 U317 ( .A(my_FIR_filter_firBlock_left_firStep[223]), .Y(n302));
   BUFX2 U318 ( .A(inData_in[3]), .Y(n303));
   BUFX2 U319 ( .A(inData_in[5]), .Y(n304));
   BUFX2 U320 ( .A(my_FIR_filter_firBlock_left_multProducts[115]), .Y(n305));
   BUFX2 U321 ( .A(my_FIR_filter_firBlock_left_multProducts[114]), .Y(n306));
   BUFX2 U322 ( .A(my_FIR_filter_firBlock_left_multProducts[113]), .Y(n307));
   BUFX2 U323 ( .A(my_FIR_filter_firBlock_left_multProducts[112]), .Y(n308));
   BUFX2 U324 ( .A(my_FIR_filter_firBlock_left_multProducts[107]), .Y(n309));
   BUFX2 U325 ( .A(my_FIR_filter_firBlock_left_multProducts[106]), .Y(n310));
   BUFX2 U326 ( .A(my_FIR_filter_firBlock_left_multProducts[105]), .Y(n311));
   BUFX2 U327 ( .A(my_FIR_filter_firBlock_left_multProducts[104]), .Y(n312));
   BUFX2 U328 ( .A(my_FIR_filter_firBlock_left_multProducts[99]), .Y(n313));
   BUFX2 U329 ( .A(my_FIR_filter_firBlock_left_multProducts[98]), .Y(n314));
   BUFX2 U330 ( .A(my_FIR_filter_firBlock_left_multProducts[97]), .Y(n315));
   BUFX2 U331 ( .A(my_FIR_filter_firBlock_left_multProducts[96]), .Y(n316));
   BUFX2 U332 ( .A(my_FIR_filter_firBlock_left_multProducts[91]), .Y(n317));
   BUFX2 U333 ( .A(leftOut[31]), .Y(n318));
   BUFX2 U334 ( .A(leftOut[30]), .Y(n319));
   BUFX2 U335 ( .A(leftOut[26]), .Y(n320));
   BUFX2 U336 ( .A(leftOut[25]), .Y(n321));
   BUFX2 U337 ( .A(leftOut[24]), .Y(n322));
   BUFX2 U338 ( .A(leftOut[23]), .Y(n323));
   BUFX2 U339 ( .A(leftOut[22]), .Y(n324));
   BUFX2 U340 ( .A(leftOut[21]), .Y(n325));
   BUFX2 U341 ( .A(leftOut[20]), .Y(n326));
   BUFX2 U342 ( .A(leftOut[19]), .Y(n327));
   BUFX2 U343 ( .A(leftOut[18]), .Y(n328));
   BUFX2 U344 ( .A(leftOut[17]), .Y(n329));
   BUFX2 U345 ( .A(leftOut[16]), .Y(n330));
   BUFX2 U346 ( .A(leftOut[15]), .Y(n331));
   BUFX2 U347 ( .A(leftOut[14]), .Y(n332));
   BUFX2 U348 ( .A(leftOut[13]), .Y(n333));
   BUFX2 U349 ( .A(leftOut[12]), .Y(n334));
   BUFX2 U350 ( .A(leftOut[11]), .Y(n335));
   BUFX2 U351 ( .A(leftOut[10]), .Y(n336));
   BUFX2 U352 ( .A(leftOut[9]), .Y(n337));
   BUFX2 U353 ( .A(leftOut[8]), .Y(n338));
   BUFX2 U354 ( .A(leftOut[7]), .Y(n339));
   BUFX2 U355 ( .A(leftOut[6]), .Y(n340));
   BUFX2 U356 ( .A(leftOut[5]), .Y(n341));
   BUFX2 U357 ( .A(leftOut[4]), .Y(n342));
   BUFX2 U358 ( .A(leftOut[3]), .Y(n343));
   BUFX2 U359 ( .A(leftOut[2]), .Y(n344));
   BUFX2 U360 ( .A(my_FIR_filter_firBlock_left_firStep[65]), .Y(n345));
   BUFX2 U361 ( .A(my_FIR_filter_firBlock_left_firStep[66]), .Y(n346));
   BUFX2 U362 ( .A(my_FIR_filter_firBlock_left_firStep[67]), .Y(n347));
   BUFX2 U363 ( .A(my_FIR_filter_firBlock_left_firStep[68]), .Y(n348));
   BUFX2 U364 ( .A(my_FIR_filter_firBlock_left_firStep[69]), .Y(n349));
   BUFX2 U365 ( .A(my_FIR_filter_firBlock_left_firStep[70]), .Y(n350));
   BUFX2 U366 ( .A(my_FIR_filter_firBlock_left_firStep[71]), .Y(n351));
   BUFX2 U367 ( .A(my_FIR_filter_firBlock_left_firStep[72]), .Y(n352));
   BUFX2 U368 ( .A(my_FIR_filter_firBlock_left_firStep[73]), .Y(n353));
   BUFX2 U369 ( .A(my_FIR_filter_firBlock_left_firStep[74]), .Y(n354));
   BUFX2 U370 ( .A(my_FIR_filter_firBlock_left_firStep[75]), .Y(n355));
   BUFX2 U371 ( .A(my_FIR_filter_firBlock_left_firStep[76]), .Y(n356));
   BUFX2 U372 ( .A(my_FIR_filter_firBlock_left_firStep[77]), .Y(n357));
   BUFX2 U373 ( .A(my_FIR_filter_firBlock_left_firStep[78]), .Y(n358));
   BUFX2 U374 ( .A(my_FIR_filter_firBlock_left_firStep[79]), .Y(n359));
   BUFX2 U375 ( .A(my_FIR_filter_firBlock_left_firStep[80]), .Y(n360));
   BUFX2 U376 ( .A(my_FIR_filter_firBlock_left_firStep[81]), .Y(n361));
   BUFX2 U377 ( .A(my_FIR_filter_firBlock_left_firStep[82]), .Y(n362));
   BUFX2 U378 ( .A(my_FIR_filter_firBlock_left_firStep[83]), .Y(n363));
   BUFX2 U379 ( .A(my_FIR_filter_firBlock_left_firStep[84]), .Y(n364));
   BUFX2 U380 ( .A(my_FIR_filter_firBlock_left_firStep[85]), .Y(n365));
   BUFX2 U381 ( .A(my_FIR_filter_firBlock_left_firStep[86]), .Y(n366));
   BUFX2 U382 ( .A(my_FIR_filter_firBlock_left_firStep[87]), .Y(n367));
   BUFX2 U383 ( .A(my_FIR_filter_firBlock_left_firStep[88]), .Y(n368));
   BUFX2 U384 ( .A(my_FIR_filter_firBlock_left_firStep[89]), .Y(n369));
   BUFX2 U385 ( .A(my_FIR_filter_firBlock_left_firStep[90]), .Y(n370));
   BUFX2 U386 ( .A(my_FIR_filter_firBlock_left_firStep[91]), .Y(n371));
   BUFX2 U387 ( .A(my_FIR_filter_firBlock_left_firStep[92]), .Y(n372));
   BUFX2 U388 ( .A(my_FIR_filter_firBlock_left_firStep[129]), .Y(n373));
   BUFX2 U389 ( .A(my_FIR_filter_firBlock_left_firStep[130]), .Y(n374));
   BUFX2 U390 ( .A(my_FIR_filter_firBlock_left_firStep[131]), .Y(n375));
   BUFX2 U391 ( .A(my_FIR_filter_firBlock_left_firStep[132]), .Y(n376));
   BUFX2 U392 ( .A(my_FIR_filter_firBlock_left_firStep[133]), .Y(n377));
   BUFX2 U393 ( .A(my_FIR_filter_firBlock_left_firStep[134]), .Y(n378));
   BUFX2 U394 ( .A(my_FIR_filter_firBlock_left_firStep[135]), .Y(n379));
   BUFX2 U395 ( .A(my_FIR_filter_firBlock_left_firStep[136]), .Y(n380));
   BUFX2 U396 ( .A(my_FIR_filter_firBlock_left_firStep[137]), .Y(n381));
   BUFX2 U397 ( .A(my_FIR_filter_firBlock_left_firStep[138]), .Y(n382));
   BUFX2 U398 ( .A(my_FIR_filter_firBlock_left_firStep[139]), .Y(n383));
   BUFX2 U399 ( .A(my_FIR_filter_firBlock_left_firStep[140]), .Y(n384));
   BUFX2 U400 ( .A(my_FIR_filter_firBlock_left_firStep[141]), .Y(n385));
   BUFX2 U401 ( .A(my_FIR_filter_firBlock_left_firStep[142]), .Y(n386));
   BUFX2 U402 ( .A(my_FIR_filter_firBlock_left_firStep[143]), .Y(n387));
   BUFX2 U403 ( .A(my_FIR_filter_firBlock_left_firStep[144]), .Y(n388));
   BUFX2 U404 ( .A(my_FIR_filter_firBlock_left_firStep[145]), .Y(n389));
   BUFX2 U405 ( .A(my_FIR_filter_firBlock_left_firStep[146]), .Y(n390));
   BUFX2 U406 ( .A(my_FIR_filter_firBlock_left_firStep[147]), .Y(n391));
   BUFX2 U407 ( .A(my_FIR_filter_firBlock_left_firStep[148]), .Y(n392));
   BUFX2 U408 ( .A(my_FIR_filter_firBlock_left_firStep[149]), .Y(n393));
   BUFX2 U409 ( .A(my_FIR_filter_firBlock_left_firStep[150]), .Y(n394));
   BUFX2 U410 ( .A(my_FIR_filter_firBlock_left_firStep[151]), .Y(n395));
   BUFX2 U411 ( .A(my_FIR_filter_firBlock_left_firStep[152]), .Y(n396));
   BUFX2 U412 ( .A(my_FIR_filter_firBlock_left_firStep[153]), .Y(n397));
   BUFX2 U413 ( .A(my_FIR_filter_firBlock_left_firStep[154]), .Y(n398));
   BUFX2 U414 ( .A(my_FIR_filter_firBlock_left_firStep[155]), .Y(n399));
   BUFX2 U415 ( .A(my_FIR_filter_firBlock_left_firStep[156]), .Y(n400));
   BUFX2 U416 ( .A(my_FIR_filter_firBlock_left_firStep[157]), .Y(n401));
   BUFX2 U417 ( .A(my_FIR_filter_firBlock_left_firStep[190]), .Y(n402));
   BUFX2 U418 ( .A(my_FIR_filter_firBlock_left_firStep[193]), .Y(n403));
   BUFX2 U419 ( .A(my_FIR_filter_firBlock_left_firStep[194]), .Y(n404));
   BUFX2 U420 ( .A(my_FIR_filter_firBlock_left_firStep[195]), .Y(n405));
   BUFX2 U421 ( .A(my_FIR_filter_firBlock_left_firStep[196]), .Y(n406));
   BUFX2 U422 ( .A(my_FIR_filter_firBlock_left_firStep[197]), .Y(n407));
   BUFX2 U423 ( .A(my_FIR_filter_firBlock_left_firStep[198]), .Y(n408));
   BUFX2 U424 ( .A(my_FIR_filter_firBlock_left_firStep[199]), .Y(n409));
   BUFX2 U425 ( .A(my_FIR_filter_firBlock_left_firStep[200]), .Y(n410));
   BUFX2 U426 ( .A(my_FIR_filter_firBlock_left_firStep[201]), .Y(n411));
   BUFX2 U427 ( .A(my_FIR_filter_firBlock_left_firStep[202]), .Y(n412));
   BUFX2 U428 ( .A(my_FIR_filter_firBlock_left_firStep[203]), .Y(n413));
   BUFX2 U429 ( .A(my_FIR_filter_firBlock_left_firStep[204]), .Y(n414));
   BUFX2 U430 ( .A(my_FIR_filter_firBlock_left_firStep[205]), .Y(n415));
   BUFX2 U431 ( .A(my_FIR_filter_firBlock_left_firStep[206]), .Y(n416));
   BUFX2 U432 ( .A(my_FIR_filter_firBlock_left_firStep[207]), .Y(n417));
   BUFX2 U433 ( .A(my_FIR_filter_firBlock_left_firStep[208]), .Y(n418));
   BUFX2 U434 ( .A(my_FIR_filter_firBlock_left_firStep[209]), .Y(n419));
   BUFX2 U435 ( .A(my_FIR_filter_firBlock_left_firStep[210]), .Y(n420));
   BUFX2 U436 ( .A(my_FIR_filter_firBlock_left_firStep[211]), .Y(n421));
   BUFX2 U437 ( .A(my_FIR_filter_firBlock_left_firStep[212]), .Y(n422));
   BUFX2 U438 ( .A(my_FIR_filter_firBlock_left_firStep[213]), .Y(n423));
   BUFX2 U439 ( .A(my_FIR_filter_firBlock_left_firStep[214]), .Y(n424));
   BUFX2 U440 ( .A(my_FIR_filter_firBlock_left_firStep[215]), .Y(n425));
   BUFX2 U441 ( .A(my_FIR_filter_firBlock_left_firStep[216]), .Y(n426));
   BUFX2 U442 ( .A(my_FIR_filter_firBlock_left_firStep[217]), .Y(n427));
   BUFX2 U443 ( .A(my_FIR_filter_firBlock_left_firStep[218]), .Y(n428));
   BUFX2 U444 ( .A(my_FIR_filter_firBlock_left_firStep[219]), .Y(n429));
   BUFX2 U445 ( .A(my_FIR_filter_firBlock_left_firStep[220]), .Y(n430));
   BUFX2 U446 ( .A(my_FIR_filter_firBlock_left_firStep[221]), .Y(n431));
   BUFX2 U447 ( .A(my_FIR_filter_firBlock_left_firStep[257]), .Y(n432));
   BUFX2 U448 ( .A(my_FIR_filter_firBlock_left_firStep[258]), .Y(n433));
   BUFX2 U449 ( .A(my_FIR_filter_firBlock_left_firStep[259]), .Y(n434));
   BUFX2 U450 ( .A(my_FIR_filter_firBlock_left_firStep[260]), .Y(n435));
   BUFX2 U451 ( .A(my_FIR_filter_firBlock_left_firStep[261]), .Y(n436));
   BUFX2 U452 ( .A(my_FIR_filter_firBlock_left_firStep[262]), .Y(n437));
   BUFX2 U453 ( .A(my_FIR_filter_firBlock_left_firStep[263]), .Y(n438));
   BUFX2 U454 ( .A(my_FIR_filter_firBlock_left_firStep[264]), .Y(n439));
   BUFX2 U455 ( .A(my_FIR_filter_firBlock_left_firStep[265]), .Y(n440));
   BUFX2 U456 ( .A(my_FIR_filter_firBlock_left_firStep[266]), .Y(n441));
   BUFX2 U457 ( .A(my_FIR_filter_firBlock_left_firStep[267]), .Y(n442));
   BUFX2 U458 ( .A(my_FIR_filter_firBlock_left_firStep[268]), .Y(n443));
   BUFX2 U459 ( .A(my_FIR_filter_firBlock_left_firStep[269]), .Y(n444));
   BUFX2 U460 ( .A(my_FIR_filter_firBlock_left_firStep[270]), .Y(n445));
   BUFX2 U461 ( .A(my_FIR_filter_firBlock_left_firStep[271]), .Y(n446));
   BUFX2 U462 ( .A(my_FIR_filter_firBlock_left_firStep[272]), .Y(n447));
   BUFX2 U463 ( .A(my_FIR_filter_firBlock_left_firStep[273]), .Y(n448));
   BUFX2 U464 ( .A(my_FIR_filter_firBlock_left_firStep[274]), .Y(n449));
   BUFX2 U465 ( .A(my_FIR_filter_firBlock_left_firStep[275]), .Y(n450));
   BUFX2 U466 ( .A(my_FIR_filter_firBlock_left_firStep[276]), .Y(n451));
   BUFX2 U467 ( .A(my_FIR_filter_firBlock_left_firStep[277]), .Y(n452));
   BUFX2 U468 ( .A(my_FIR_filter_firBlock_left_firStep[278]), .Y(n453));
   BUFX2 U469 ( .A(my_FIR_filter_firBlock_left_firStep[279]), .Y(n454));
   BUFX2 U470 ( .A(my_FIR_filter_firBlock_left_firStep[280]), .Y(n455));
   BUFX2 U471 ( .A(my_FIR_filter_firBlock_left_firStep[281]), .Y(n456));
   BUFX2 U472 ( .A(my_FIR_filter_firBlock_left_firStep[282]), .Y(n457));
   BUFX2 U473 ( .A(my_FIR_filter_firBlock_left_firStep[283]), .Y(n458));
   BUFX2 U474 ( .A(my_FIR_filter_firBlock_left_firStep[284]), .Y(n459));
   BUFX2 U475 ( .A(leftOut[27]), .Y(n460));
   BUFX2 U476 ( .A(leftOut[29]), .Y(n461));
   BUFX2 U477 ( .A(leftOut[28]), .Y(n462));
   BUFX2 U478 ( .A(leftOut[1]), .Y(n463));
   BUFX2 U479 ( .A(my_FIR_filter_firBlock_left_firStep[64]), .Y(n464));
   BUFX2 U480 ( .A(my_FIR_filter_firBlock_left_firStep[128]), .Y(n465));
   BUFX2 U481 ( .A(my_FIR_filter_firBlock_left_firStep[192]), .Y(n466));
   BUFX2 U482 ( .A(my_FIR_filter_firBlock_left_firStep[256]), .Y(n467));
   BUFX2 U483 ( .A(leftOut[0]), .Y(n468));
   BUFX2 U484 ( .A(my_FIR_filter_firBlock_left_firStep[63]), .Y(n469));
   BUFX2 U485 ( .A(my_FIR_filter_firBlock_left_firStep[127]), .Y(n470));
   BUFX2 U486 ( .A(my_FIR_filter_firBlock_left_firStep[191]), .Y(n471));
   BUFX2 U487 ( .A(my_FIR_filter_firBlock_left_firStep[255]), .Y(n472));
   BUFX2 U488 ( .A(inData_in[2]), .Y(n473));
   BUFX2 U489 ( .A(my_FIR_filter_firBlock_left_multProducts[111]), .Y(n474));
   BUFX2 U490 ( .A(my_FIR_filter_firBlock_left_multProducts[110]), .Y(n475));
   BUFX2 U491 ( .A(my_FIR_filter_firBlock_left_multProducts[109]), .Y(n476));
   BUFX2 U492 ( .A(my_FIR_filter_firBlock_left_multProducts[108]), .Y(n477));
   BUFX2 U493 ( .A(my_FIR_filter_firBlock_left_multProducts[103]), .Y(n478));
   BUFX2 U494 ( .A(my_FIR_filter_firBlock_left_multProducts[102]), .Y(n479));
   BUFX2 U495 ( .A(my_FIR_filter_firBlock_left_multProducts[101]), .Y(n480));
   BUFX2 U496 ( .A(my_FIR_filter_firBlock_left_multProducts[100]), .Y(n481));
   BUFX2 U497 ( .A(my_FIR_filter_firBlock_left_multProducts[95]), .Y(n482));
   BUFX2 U498 ( .A(my_FIR_filter_firBlock_left_multProducts[93]), .Y(n483));
   BUFX2 U499 ( .A(my_FIR_filter_firBlock_left_multProducts[94]), .Y(n484));
   BUFX2 U500 ( .A(my_FIR_filter_firBlock_left_multProducts[92]), .Y(n485));
   BUFX2 U501 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_134_carry[36]), .Y(n486));
   AND2X1 U502 ( .A(n603),  .B(n515), .Y(n487));
   AND2X1 U503 ( .A(n602),  .B(n487), .Y(n488));
   AND2X1 U504 ( .A(n601),  .B(n488), .Y(n489));
   AND2X1 U505 ( .A(n600),  .B(n489), .Y(n490));
   AND2X1 U506 ( .A(n599),  .B(n490), .Y(n491));
   AND2X1 U507 ( .A(n598),  .B(n491), .Y(n492));
   AND2X1 U508 ( .A(n597),  .B(n492), .Y(n493));
   AND2X1 U509 ( .A(n596),  .B(n493), .Y(n494));
   AND2X1 U510 ( .A(n595),  .B(n494), .Y(n495));
   AND2X1 U511 ( .A(n594),  .B(n495), .Y(n496));
   AND2X1 U512 ( .A(n593),  .B(n496), .Y(n497));
   AND2X1 U513 ( .A(n592),  .B(n497), .Y(n498));
   AND2X1 U514 ( .A(n591),  .B(n498), .Y(n499));
   AND2X1 U515 ( .A(n590),  .B(n499), .Y(n500));
   AND2X1 U516 ( .A(n589),  .B(n500), .Y(n501));
   AND2X1 U517 ( .A(n588),  .B(n501), .Y(n502));
   AND2X1 U518 ( .A(n587),  .B(n502), .Y(n503));
   AND2X1 U519 ( .A(n586),  .B(n503), .Y(n504));
   AND2X1 U520 ( .A(n585),  .B(n504), .Y(n505));
   AND2X1 U521 ( .A(n584),  .B(n505), .Y(n506));
   AND2X1 U522 ( .A(n583),  .B(n506), .Y(n507));
   AND2X1 U523 ( .A(n582),  .B(n507), .Y(n508));
   AND2X1 U524 ( .A(n581),  .B(n508), .Y(n509));
   AND2X1 U525 ( .A(n580),  .B(n509), .Y(n510));
   AND2X1 U526 ( .A(n579),  .B(n510), .Y(n511));
   AND2X1 U527 ( .A(n578),  .B(n511), .Y(n512));
   AND2X1 U528 ( .A(n577),  .B(n512), .Y(n513));
   AND2X1 U529 ( .A(n576),  .B(n513), .Y(n514));
   AND2X1 U530 ( .A(n604),  .B(n605), .Y(n515));
   AND2X1 U531 ( .A(n573),  .B(n572), .Y(n517));
   XOR2X1 U532 ( .A(n604),  .B(n605), .Y(puf_84_wire_1));
   XOR2X1 U533 ( .A(n603),  .B(n515), .Y(puf_85_wire_1));
   XOR2X1 U534 ( .A(n602),  .B(n487), .Y(puf_86_wire_1));
   XOR2X1 U535 ( .A(n601),  .B(n488), .Y(puf_87_wire_1));
   XOR2X1 U536 ( .A(n600),  .B(n489), .Y(puf_88_wire_1));
   XOR2X1 U537 ( .A(n599),  .B(n490), .Y(puf_89_wire_1));
   XOR2X1 U538 ( .A(n598),  .B(n491), .Y(puf_90_wire_1));
   XOR2X1 U539 ( .A(n597),  .B(n492), .Y(puf_91_wire_1));
   XOR2X1 U540 ( .A(n596),  .B(n493), .Y(puf_92_wire_1));
   XOR2X1 U541 ( .A(n595),  .B(n494), .Y(puf_93_wire_1));
   XOR2X1 U542 ( .A(n594),  .B(n495), .Y(puf_94_wire_1));
   XOR2X1 U543 ( .A(n593),  .B(n496), .Y(puf_95_wire_1));
   XOR2X1 U544 ( .A(n592),  .B(n497), .Y(puf_96_wire_1));
   XOR2X1 U545 ( .A(n591),  .B(n498), .Y(puf_97_wire_1));
   XOR2X1 U546 ( .A(n590),  .B(n499), .Y(puf_98_wire_1));
   XOR2X1 U547 ( .A(n589),  .B(n500), .Y(puf_99_wire_1));
   XOR2X1 U548 ( .A(n588),  .B(n501), .Y(puf_100_wire_1));
   XOR2X1 U549 ( .A(n587),  .B(n502), .Y(puf_101_wire_1));
   XOR2X1 U550 ( .A(n586),  .B(n503), .Y(puf_102_wire_1));
   XOR2X1 U551 ( .A(n585),  .B(n504), .Y(my_FIR_filter_firBlock_right_multProducts[20]));
   XOR2X1 U552 ( .A(n584),  .B(n505), .Y(my_FIR_filter_firBlock_right_multProducts[21]));
   XOR2X1 U553 ( .A(n583),  .B(n506), .Y(my_FIR_filter_firBlock_right_multProducts[22]));
   XOR2X1 U554 ( .A(n582),  .B(n507), .Y(my_FIR_filter_firBlock_right_multProducts[23]));
   XOR2X1 U555 ( .A(n581),  .B(n508), .Y(my_FIR_filter_firBlock_right_multProducts[24]));
   XOR2X1 U556 ( .A(n580),  .B(n509), .Y(my_FIR_filter_firBlock_right_multProducts[25]));
   XOR2X1 U557 ( .A(n579),  .B(n510), .Y(my_FIR_filter_firBlock_right_multProducts[26]));
   XOR2X1 U558 ( .A(n578),  .B(n511), .Y(my_FIR_filter_firBlock_right_multProducts[27]));
   XOR2X1 U559 ( .A(n577),  .B(n512), .Y(my_FIR_filter_firBlock_right_multProducts[28]));
   XOR2X1 U560 ( .A(n576),  .B(n513), .Y(my_FIR_filter_firBlock_right_multProducts[29]));
   XOR2X1 U561 ( .A(n575),  .B(n514), .Y(my_FIR_filter_firBlock_right_multProducts[30]));
   XOR2X1 U562 ( .A(n574),  .B(n527), .Y(my_FIR_filter_firBlock_right_multProducts[31]));
   XOR2X1 U563 ( .A(my_FIR_filter_firBlock_left_multProducts[62]),  .B(n136), .Y(puf_103_wire_1));
   XOR2X1 U564 ( .A(my_FIR_filter_firBlock_left_multProducts[33]),  .B(n472), .Y(puf_104_wire_1));
   XOR2X1 U565 ( .A(my_FIR_filter_firBlock_left_multProducts[32]),  .B(n302), .Y(puf_105_wire_1));
   XOR2X1 U566 ( .A(my_FIR_filter_firBlock_left_multProducts[0]),  .B(n471), .Y(puf_106_wire_1));
   XOR2X1 U567 ( .A(my_FIR_filter_firBlock_left_multProducts[0]),  .B(n301), .Y(puf_107_wire_1));
   XOR2X1 U568 ( .A(my_FIR_filter_firBlock_left_multProducts[32]),  .B(n470), .Y(puf_108_wire_1));
   XOR2X1 U569 ( .A(my_FIR_filter_firBlock_left_multProducts[33]),  .B(n300), .Y(puf_109_wire_1));
   XOR2X1 U570 ( .A(my_FIR_filter_firBlock_left_multProducts[62]),  .B(n469), .Y(puf_110_wire_1));
   XOR2X1 U571 ( .A(n317),  .B(n135), .Y(puf_111_wire_1));
   XOR2X1 U572 ( .A(n299),  .B(n468), .Y(outData_in[0]));
   INVX1 U573 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_138_carry[33]), .Y(n541));
   INVX1 U574 ( .A(n486), .Y(n542));
   INVX1 U575 ( .A(n305), .Y(n543));
   INVX1 U576 ( .A(n306), .Y(n544));
   INVX1 U577 ( .A(n307), .Y(n545));
   INVX1 U578 ( .A(n308), .Y(n546));
   INVX1 U579 ( .A(n474), .Y(n547));
   INVX1 U580 ( .A(n475), .Y(n548));
   INVX1 U581 ( .A(n476), .Y(n549));
   INVX1 U582 ( .A(n477), .Y(n550));
   INVX1 U583 ( .A(n309), .Y(n551));
   INVX1 U584 ( .A(n310), .Y(n552));
   INVX1 U585 ( .A(n311), .Y(n553));
   INVX1 U586 ( .A(n312), .Y(n554));
   INVX1 U587 ( .A(n478), .Y(n555));
   INVX1 U588 ( .A(n479), .Y(n556));
   INVX1 U589 ( .A(n480), .Y(n557));
   INVX1 U590 ( .A(n481), .Y(n558));
   INVX1 U591 ( .A(n313), .Y(n559));
   INVX1 U592 ( .A(n314), .Y(n560));
   INVX1 U593 ( .A(n315), .Y(n561));
   INVX1 U594 ( .A(n316), .Y(n562));
   INVX1 U595 ( .A(n482), .Y(n563));
   INVX1 U596 ( .A(n484), .Y(n564));
   INVX1 U597 ( .A(n483), .Y(n565));
   INVX1 U598 ( .A(n485), .Y(n566));
   INVX1 U599 ( .A(n317), .Y(n567));
   INVX1 U600 ( .A(n103), .Y(n573));
   INVX1 U601 ( .A(outData_in[31]), .Y(n574));
   INVX1 U602 ( .A(outData_in[30]), .Y(n575));
   INVX1 U603 ( .A(outData_in[29]), .Y(n576));
   INVX1 U604 ( .A(outData_in[28]), .Y(n577));
   INVX1 U605 ( .A(outData_in[27]), .Y(n578));
   INVX1 U606 ( .A(outData_in[26]), .Y(n579));
   INVX1 U607 ( .A(outData_in[25]), .Y(n580));
   INVX1 U608 ( .A(outData_in[24]), .Y(n581));
   INVX1 U609 ( .A(outData_in[23]), .Y(n582));
   INVX1 U610 ( .A(outData_in[22]), .Y(n583));
   INVX1 U611 ( .A(outData_in[21]), .Y(n584));
   INVX1 U612 ( .A(outData_in[20]), .Y(n585));
   INVX1 U613 ( .A(outData_in[19]), .Y(n586));
   INVX1 U614 ( .A(outData_in[18]), .Y(n587));
   INVX1 U615 ( .A(outData_in[17]), .Y(n588));
   INVX1 U616 ( .A(outData_in[16]), .Y(n589));
   INVX1 U617 ( .A(outData_in[15]), .Y(n590));
   INVX1 U618 ( .A(outData_in[14]), .Y(n591));
   INVX1 U619 ( .A(outData_in[13]), .Y(n592));
   INVX1 U620 ( .A(outData_in[12]), .Y(n593));
   INVX1 U621 ( .A(outData_in[11]), .Y(n594));
   INVX1 U622 ( .A(outData_in[10]), .Y(n595));
   INVX1 U623 ( .A(outData_in[9]), .Y(n596));
   INVX1 U624 ( .A(outData_in[8]), .Y(n597));
   INVX1 U625 ( .A(outData_in[7]), .Y(n598));
   INVX1 U626 ( .A(outData_in[6]), .Y(n599));
   INVX1 U627 ( .A(outData_in[5]), .Y(n600));
   INVX1 U628 ( .A(outData_in[4]), .Y(n601));
   INVX1 U629 ( .A(outData_in[3]), .Y(n602));
   INVX1 U630 ( .A(outData_in[2]), .Y(n603));
   INVX1 U631 ( .A(outData_in[1]), .Y(n604));
   INVX1 U632 ( .A(outData_in[0]), .Y(n605));
   OAI21X1 U633 ( .A(n485),  .B(n66),  .C(n528), .Y(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_sub_135_carry[8]));
   OAI21X1 U634 ( .A(n529),  .B(n103),  .C(n99), .Y(n528));
   AOI21X1 U635 ( .A(n485),  .B(n66),  .C(n317), .Y(n530));
   NOR3X1 U636 ( .A(n100),  .B(n473),  .C(n137), .Y(n529));
   NAND3X1 U637 ( .A(n569),  .B(n568),  .C(n570), .Y(n531));
   INVX1 U638 ( .A(n304), .Y(n568));
   INVX1 U639 ( .A(n138), .Y(n569));
   OAI21X1 U640 ( .A(n570),  .B(n532),  .C(n533), .Y(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_add_131_carry[7]));
   OAI21X1 U641 ( .A(n303),  .B(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_12_),  .C(n534), .Y(n533));
   OAI21X1 U642 ( .A(n571),  .B(n535),  .C(n536), .Y(n534));
   OAI21X1 U643 ( .A(n473),  .B(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_11_),  .C(n537), .Y(n536));
   OAI21X1 U644 ( .A(n572),  .B(n538),  .C(n101), .Y(n537));
   NAND3X1 U645 ( .A(n102),  .B(n103),  .C(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_9_), .Y(n539));
   INVX1 U646 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_10_), .Y(n538));
   INVX1 U647 ( .A(n137), .Y(n572));
   INVX1 U648 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_11_), .Y(n535));
   INVX1 U649 ( .A(n473), .Y(n571));
   INVX1 U650 ( .A(my_FIR_filter_firBlock_left_my_FIR_filter_firBlock_left_MultiplyBlock_w192_12_), .Y(n532));
   INVX1 U651 ( .A(n303), .Y(n570));
   INVX1 puf_0_instance_0 ( .A(puf_0_wire_1), .Y(puf_0_wire_0));
   MUX2X1 puf_0_instance_1 ( .A(puf_0_wire_0),  .B(outData[31]),  .S(sel), .Y(puf_0_wire_2));
   INVX1 puf_0_instance_2 ( .A(puf_0_wire_2), .Y(puf_0_wire_5));
   INVX1 puf_0_instance_3 ( .A(puf_0_wire_5), .Y(puf_0_wire_6));
   MUX2X1 puf_0_instance_4 ( .A(puf_0_wire_0),  .B(puf_0_wire_6),  .S(sel), .Y(puf_0_wire_7));
   INVX1 puf_0_instance_5 ( .A(puf_0_wire_7), .Y(puf_0_wire_8));
   INVX1 puf_0_instance_6 ( .A(puf_0_wire_8), .Y(outData[31]));
   BUFX2 puf_out_instance_0 ( .A(outData[31]), .Y(pufout[0]));
   INVX1 puf_1_instance_0 ( .A(puf_1_wire_1), .Y(puf_1_wire_0));
   MUX2X1 puf_1_instance_1 ( .A(puf_1_wire_0),  .B(outData[30]),  .S(sel), .Y(puf_1_wire_2));
   INVX1 puf_1_instance_2 ( .A(puf_1_wire_2), .Y(puf_1_wire_5));
   INVX1 puf_1_instance_3 ( .A(puf_1_wire_5), .Y(puf_1_wire_6));
   MUX2X1 puf_1_instance_4 ( .A(puf_1_wire_0),  .B(puf_1_wire_6),  .S(sel), .Y(puf_1_wire_7));
   INVX1 puf_1_instance_5 ( .A(puf_1_wire_7), .Y(puf_1_wire_8));
   INVX1 puf_1_instance_6 ( .A(puf_1_wire_8), .Y(outData[30]));
   BUFX2 puf_out_instance_1 ( .A(outData[30]), .Y(pufout[1]));
   INVX1 puf_2_instance_0 ( .A(puf_2_wire_1), .Y(puf_2_wire_0));
   MUX2X1 puf_2_instance_1 ( .A(puf_2_wire_0),  .B(outData[29]),  .S(sel), .Y(puf_2_wire_2));
   INVX1 puf_2_instance_2 ( .A(puf_2_wire_2), .Y(puf_2_wire_5));
   INVX1 puf_2_instance_3 ( .A(puf_2_wire_5), .Y(puf_2_wire_6));
   MUX2X1 puf_2_instance_4 ( .A(puf_2_wire_0),  .B(puf_2_wire_6),  .S(sel), .Y(puf_2_wire_7));
   INVX1 puf_2_instance_5 ( .A(puf_2_wire_7), .Y(puf_2_wire_8));
   INVX1 puf_2_instance_6 ( .A(puf_2_wire_8), .Y(outData[29]));
   BUFX2 puf_out_instance_2 ( .A(outData[29]), .Y(pufout[2]));
   INVX1 puf_3_instance_0 ( .A(puf_3_wire_1), .Y(puf_3_wire_0));
   MUX2X1 puf_3_instance_1 ( .A(puf_3_wire_0),  .B(outData[28]),  .S(sel), .Y(puf_3_wire_2));
   INVX1 puf_3_instance_2 ( .A(puf_3_wire_2), .Y(puf_3_wire_5));
   INVX1 puf_3_instance_3 ( .A(puf_3_wire_5), .Y(puf_3_wire_6));
   MUX2X1 puf_3_instance_4 ( .A(puf_3_wire_0),  .B(puf_3_wire_6),  .S(sel), .Y(puf_3_wire_7));
   INVX1 puf_3_instance_5 ( .A(puf_3_wire_7), .Y(puf_3_wire_8));
   INVX1 puf_3_instance_6 ( .A(puf_3_wire_8), .Y(outData[28]));
   BUFX2 puf_out_instance_3 ( .A(outData[28]), .Y(pufout[3]));
   INVX1 puf_4_instance_0 ( .A(puf_4_wire_1), .Y(puf_4_wire_0));
   MUX2X1 puf_4_instance_1 ( .A(puf_4_wire_0),  .B(outData[27]),  .S(sel), .Y(puf_4_wire_2));
   INVX1 puf_4_instance_2 ( .A(puf_4_wire_2), .Y(puf_4_wire_5));
   INVX1 puf_4_instance_3 ( .A(puf_4_wire_5), .Y(puf_4_wire_6));
   MUX2X1 puf_4_instance_4 ( .A(puf_4_wire_0),  .B(puf_4_wire_6),  .S(sel), .Y(puf_4_wire_7));
   INVX1 puf_4_instance_5 ( .A(puf_4_wire_7), .Y(puf_4_wire_8));
   INVX1 puf_4_instance_6 ( .A(puf_4_wire_8), .Y(outData[27]));
   BUFX2 puf_out_instance_4 ( .A(outData[27]), .Y(pufout[4]));
   INVX1 puf_5_instance_0 ( .A(puf_5_wire_1), .Y(puf_5_wire_0));
   MUX2X1 puf_5_instance_1 ( .A(puf_5_wire_0),  .B(outData[26]),  .S(sel), .Y(puf_5_wire_2));
   INVX1 puf_5_instance_2 ( .A(puf_5_wire_2), .Y(puf_5_wire_5));
   INVX1 puf_5_instance_3 ( .A(puf_5_wire_5), .Y(puf_5_wire_6));
   MUX2X1 puf_5_instance_4 ( .A(puf_5_wire_0),  .B(puf_5_wire_6),  .S(sel), .Y(puf_5_wire_7));
   INVX1 puf_5_instance_5 ( .A(puf_5_wire_7), .Y(puf_5_wire_8));
   INVX1 puf_5_instance_6 ( .A(puf_5_wire_8), .Y(outData[26]));
   BUFX2 puf_out_instance_5 ( .A(outData[26]), .Y(pufout[5]));
   INVX1 puf_6_instance_0 ( .A(puf_6_wire_1), .Y(puf_6_wire_0));
   MUX2X1 puf_6_instance_1 ( .A(puf_6_wire_0),  .B(outData[25]),  .S(sel), .Y(puf_6_wire_2));
   INVX1 puf_6_instance_2 ( .A(puf_6_wire_2), .Y(puf_6_wire_5));
   INVX1 puf_6_instance_3 ( .A(puf_6_wire_5), .Y(puf_6_wire_6));
   MUX2X1 puf_6_instance_4 ( .A(puf_6_wire_0),  .B(puf_6_wire_6),  .S(sel), .Y(puf_6_wire_7));
   INVX1 puf_6_instance_5 ( .A(puf_6_wire_7), .Y(puf_6_wire_8));
   INVX1 puf_6_instance_6 ( .A(puf_6_wire_8), .Y(outData[25]));
   BUFX2 puf_out_instance_6 ( .A(outData[25]), .Y(pufout[6]));
   INVX1 puf_7_instance_0 ( .A(puf_7_wire_1), .Y(puf_7_wire_0));
   MUX2X1 puf_7_instance_1 ( .A(puf_7_wire_0),  .B(outData[24]),  .S(sel), .Y(puf_7_wire_2));
   INVX1 puf_7_instance_2 ( .A(puf_7_wire_2), .Y(puf_7_wire_5));
   INVX1 puf_7_instance_3 ( .A(puf_7_wire_5), .Y(puf_7_wire_6));
   MUX2X1 puf_7_instance_4 ( .A(puf_7_wire_0),  .B(puf_7_wire_6),  .S(sel), .Y(puf_7_wire_7));
   INVX1 puf_7_instance_5 ( .A(puf_7_wire_7), .Y(puf_7_wire_8));
   INVX1 puf_7_instance_6 ( .A(puf_7_wire_8), .Y(outData[24]));
   BUFX2 puf_out_instance_7 ( .A(outData[24]), .Y(pufout[7]));
   INVX1 puf_8_instance_0 ( .A(puf_8_wire_1), .Y(puf_8_wire_0));
   MUX2X1 puf_8_instance_1 ( .A(puf_8_wire_0),  .B(outData[23]),  .S(sel), .Y(puf_8_wire_2));
   INVX1 puf_8_instance_2 ( .A(puf_8_wire_2), .Y(puf_8_wire_5));
   INVX1 puf_8_instance_3 ( .A(puf_8_wire_5), .Y(puf_8_wire_6));
   MUX2X1 puf_8_instance_4 ( .A(puf_8_wire_0),  .B(puf_8_wire_6),  .S(sel), .Y(puf_8_wire_7));
   INVX1 puf_8_instance_5 ( .A(puf_8_wire_7), .Y(puf_8_wire_8));
   INVX1 puf_8_instance_6 ( .A(puf_8_wire_8), .Y(outData[23]));
   BUFX2 puf_out_instance_8 ( .A(outData[23]), .Y(pufout[8]));
   INVX1 puf_9_instance_0 ( .A(puf_9_wire_1), .Y(puf_9_wire_0));
   MUX2X1 puf_9_instance_1 ( .A(puf_9_wire_0),  .B(outData[22]),  .S(sel), .Y(puf_9_wire_2));
   INVX1 puf_9_instance_2 ( .A(puf_9_wire_2), .Y(puf_9_wire_5));
   INVX1 puf_9_instance_3 ( .A(puf_9_wire_5), .Y(puf_9_wire_6));
   MUX2X1 puf_9_instance_4 ( .A(puf_9_wire_0),  .B(puf_9_wire_6),  .S(sel), .Y(puf_9_wire_7));
   INVX1 puf_9_instance_5 ( .A(puf_9_wire_7), .Y(puf_9_wire_8));
   INVX1 puf_9_instance_6 ( .A(puf_9_wire_8), .Y(outData[22]));
   BUFX2 puf_out_instance_9 ( .A(outData[22]), .Y(pufout[9]));
   INVX1 puf_10_instance_0 ( .A(puf_10_wire_1), .Y(puf_10_wire_0));
   MUX2X1 puf_10_instance_1 ( .A(puf_10_wire_0),  .B(outData[21]),  .S(sel), .Y(puf_10_wire_2));
   INVX1 puf_10_instance_2 ( .A(puf_10_wire_2), .Y(puf_10_wire_5));
   INVX1 puf_10_instance_3 ( .A(puf_10_wire_5), .Y(puf_10_wire_6));
   MUX2X1 puf_10_instance_4 ( .A(puf_10_wire_0),  .B(puf_10_wire_6),  .S(sel), .Y(puf_10_wire_7));
   INVX1 puf_10_instance_5 ( .A(puf_10_wire_7), .Y(puf_10_wire_8));
   INVX1 puf_10_instance_6 ( .A(puf_10_wire_8), .Y(outData[21]));
   BUFX2 puf_out_instance_10 ( .A(outData[21]), .Y(pufout[10]));
   INVX1 puf_11_instance_0 ( .A(puf_11_wire_1), .Y(puf_11_wire_0));
   MUX2X1 puf_11_instance_1 ( .A(puf_11_wire_0),  .B(outData[20]),  .S(sel), .Y(puf_11_wire_2));
   INVX1 puf_11_instance_2 ( .A(puf_11_wire_2), .Y(puf_11_wire_5));
   INVX1 puf_11_instance_3 ( .A(puf_11_wire_5), .Y(puf_11_wire_6));
   MUX2X1 puf_11_instance_4 ( .A(puf_11_wire_0),  .B(puf_11_wire_6),  .S(sel), .Y(puf_11_wire_7));
   INVX1 puf_11_instance_5 ( .A(puf_11_wire_7), .Y(puf_11_wire_8));
   INVX1 puf_11_instance_6 ( .A(puf_11_wire_8), .Y(outData[20]));
   BUFX2 puf_out_instance_11 ( .A(outData[20]), .Y(pufout[11]));
   INVX1 puf_12_instance_0 ( .A(puf_12_wire_1), .Y(puf_12_wire_0));
   MUX2X1 puf_12_instance_1 ( .A(puf_12_wire_0),  .B(outData[19]),  .S(sel), .Y(puf_12_wire_2));
   INVX1 puf_12_instance_2 ( .A(puf_12_wire_2), .Y(puf_12_wire_5));
   INVX1 puf_12_instance_3 ( .A(puf_12_wire_5), .Y(puf_12_wire_6));
   MUX2X1 puf_12_instance_4 ( .A(puf_12_wire_0),  .B(puf_12_wire_6),  .S(sel), .Y(puf_12_wire_7));
   INVX1 puf_12_instance_5 ( .A(puf_12_wire_7), .Y(puf_12_wire_8));
   INVX1 puf_12_instance_6 ( .A(puf_12_wire_8), .Y(outData[19]));
   BUFX2 puf_out_instance_12 ( .A(outData[19]), .Y(pufout[12]));
   INVX1 puf_13_instance_0 ( .A(puf_13_wire_1), .Y(puf_13_wire_0));
   MUX2X1 puf_13_instance_1 ( .A(puf_13_wire_0),  .B(outData[18]),  .S(sel), .Y(puf_13_wire_2));
   INVX1 puf_13_instance_2 ( .A(puf_13_wire_2), .Y(puf_13_wire_5));
   INVX1 puf_13_instance_3 ( .A(puf_13_wire_5), .Y(puf_13_wire_6));
   MUX2X1 puf_13_instance_4 ( .A(puf_13_wire_0),  .B(puf_13_wire_6),  .S(sel), .Y(puf_13_wire_7));
   INVX1 puf_13_instance_5 ( .A(puf_13_wire_7), .Y(puf_13_wire_8));
   INVX1 puf_13_instance_6 ( .A(puf_13_wire_8), .Y(outData[18]));
   BUFX2 puf_out_instance_13 ( .A(outData[18]), .Y(pufout[13]));
   INVX1 puf_14_instance_0 ( .A(puf_14_wire_1), .Y(puf_14_wire_0));
   MUX2X1 puf_14_instance_1 ( .A(puf_14_wire_0),  .B(outData[17]),  .S(sel), .Y(puf_14_wire_2));
   INVX1 puf_14_instance_2 ( .A(puf_14_wire_2), .Y(puf_14_wire_5));
   INVX1 puf_14_instance_3 ( .A(puf_14_wire_5), .Y(puf_14_wire_6));
   MUX2X1 puf_14_instance_4 ( .A(puf_14_wire_0),  .B(puf_14_wire_6),  .S(sel), .Y(puf_14_wire_7));
   INVX1 puf_14_instance_5 ( .A(puf_14_wire_7), .Y(puf_14_wire_8));
   INVX1 puf_14_instance_6 ( .A(puf_14_wire_8), .Y(outData[17]));
   BUFX2 puf_out_instance_14 ( .A(outData[17]), .Y(pufout[14]));
   INVX1 puf_15_instance_0 ( .A(puf_15_wire_1), .Y(puf_15_wire_0));
   MUX2X1 puf_15_instance_1 ( .A(puf_15_wire_0),  .B(outData[16]),  .S(sel), .Y(puf_15_wire_2));
   INVX1 puf_15_instance_2 ( .A(puf_15_wire_2), .Y(puf_15_wire_5));
   INVX1 puf_15_instance_3 ( .A(puf_15_wire_5), .Y(puf_15_wire_6));
   MUX2X1 puf_15_instance_4 ( .A(puf_15_wire_0),  .B(puf_15_wire_6),  .S(sel), .Y(puf_15_wire_7));
   INVX1 puf_15_instance_5 ( .A(puf_15_wire_7), .Y(puf_15_wire_8));
   INVX1 puf_15_instance_6 ( .A(puf_15_wire_8), .Y(outData[16]));
   BUFX2 puf_out_instance_15 ( .A(outData[16]), .Y(pufout[15]));
   INVX1 puf_16_instance_0 ( .A(puf_16_wire_1), .Y(puf_16_wire_0));
   MUX2X1 puf_16_instance_1 ( .A(puf_16_wire_0),  .B(outData[15]),  .S(sel), .Y(puf_16_wire_2));
   INVX1 puf_16_instance_2 ( .A(puf_16_wire_2), .Y(puf_16_wire_5));
   INVX1 puf_16_instance_3 ( .A(puf_16_wire_5), .Y(puf_16_wire_6));
   MUX2X1 puf_16_instance_4 ( .A(puf_16_wire_0),  .B(puf_16_wire_6),  .S(sel), .Y(puf_16_wire_7));
   INVX1 puf_16_instance_5 ( .A(puf_16_wire_7), .Y(puf_16_wire_8));
   INVX1 puf_16_instance_6 ( .A(puf_16_wire_8), .Y(outData[15]));
   BUFX2 puf_out_instance_16 ( .A(outData[15]), .Y(pufout[16]));
   INVX1 puf_17_instance_0 ( .A(puf_17_wire_1), .Y(puf_17_wire_0));
   MUX2X1 puf_17_instance_1 ( .A(puf_17_wire_0),  .B(outData[14]),  .S(sel), .Y(puf_17_wire_2));
   INVX1 puf_17_instance_2 ( .A(puf_17_wire_2), .Y(puf_17_wire_5));
   INVX1 puf_17_instance_3 ( .A(puf_17_wire_5), .Y(puf_17_wire_6));
   MUX2X1 puf_17_instance_4 ( .A(puf_17_wire_0),  .B(puf_17_wire_6),  .S(sel), .Y(puf_17_wire_7));
   INVX1 puf_17_instance_5 ( .A(puf_17_wire_7), .Y(puf_17_wire_8));
   INVX1 puf_17_instance_6 ( .A(puf_17_wire_8), .Y(outData[14]));
   BUFX2 puf_out_instance_17 ( .A(outData[14]), .Y(pufout[17]));
   INVX1 puf_18_instance_0 ( .A(puf_18_wire_1), .Y(puf_18_wire_0));
   MUX2X1 puf_18_instance_1 ( .A(puf_18_wire_0),  .B(outData[13]),  .S(sel), .Y(puf_18_wire_2));
   INVX1 puf_18_instance_2 ( .A(puf_18_wire_2), .Y(puf_18_wire_5));
   INVX1 puf_18_instance_3 ( .A(puf_18_wire_5), .Y(puf_18_wire_6));
   MUX2X1 puf_18_instance_4 ( .A(puf_18_wire_0),  .B(puf_18_wire_6),  .S(sel), .Y(puf_18_wire_7));
   INVX1 puf_18_instance_5 ( .A(puf_18_wire_7), .Y(puf_18_wire_8));
   INVX1 puf_18_instance_6 ( .A(puf_18_wire_8), .Y(outData[13]));
   BUFX2 puf_out_instance_18 ( .A(outData[13]), .Y(pufout[18]));
   INVX1 puf_19_instance_0 ( .A(puf_19_wire_1), .Y(puf_19_wire_0));
   MUX2X1 puf_19_instance_1 ( .A(puf_19_wire_0),  .B(outData[12]),  .S(sel), .Y(puf_19_wire_2));
   INVX1 puf_19_instance_2 ( .A(puf_19_wire_2), .Y(puf_19_wire_5));
   INVX1 puf_19_instance_3 ( .A(puf_19_wire_5), .Y(puf_19_wire_6));
   MUX2X1 puf_19_instance_4 ( .A(puf_19_wire_0),  .B(puf_19_wire_6),  .S(sel), .Y(puf_19_wire_7));
   INVX1 puf_19_instance_5 ( .A(puf_19_wire_7), .Y(puf_19_wire_8));
   INVX1 puf_19_instance_6 ( .A(puf_19_wire_8), .Y(outData[12]));
   BUFX2 puf_out_instance_19 ( .A(outData[12]), .Y(pufout[19]));
   INVX1 puf_20_instance_0 ( .A(puf_20_wire_1), .Y(puf_20_wire_0));
   MUX2X1 puf_20_instance_1 ( .A(puf_20_wire_0),  .B(outData[11]),  .S(sel), .Y(puf_20_wire_2));
   INVX1 puf_20_instance_2 ( .A(puf_20_wire_2), .Y(puf_20_wire_5));
   INVX1 puf_20_instance_3 ( .A(puf_20_wire_5), .Y(puf_20_wire_6));
   MUX2X1 puf_20_instance_4 ( .A(puf_20_wire_0),  .B(puf_20_wire_6),  .S(sel), .Y(puf_20_wire_7));
   INVX1 puf_20_instance_5 ( .A(puf_20_wire_7), .Y(puf_20_wire_8));
   INVX1 puf_20_instance_6 ( .A(puf_20_wire_8), .Y(outData[11]));
   BUFX2 puf_out_instance_20 ( .A(outData[11]), .Y(pufout[20]));
   INVX1 puf_21_instance_0 ( .A(puf_21_wire_1), .Y(puf_21_wire_0));
   MUX2X1 puf_21_instance_1 ( .A(puf_21_wire_0),  .B(outData[10]),  .S(sel), .Y(puf_21_wire_2));
   INVX1 puf_21_instance_2 ( .A(puf_21_wire_2), .Y(puf_21_wire_5));
   INVX1 puf_21_instance_3 ( .A(puf_21_wire_5), .Y(puf_21_wire_6));
   MUX2X1 puf_21_instance_4 ( .A(puf_21_wire_0),  .B(puf_21_wire_6),  .S(sel), .Y(puf_21_wire_7));
   INVX1 puf_21_instance_5 ( .A(puf_21_wire_7), .Y(puf_21_wire_8));
   INVX1 puf_21_instance_6 ( .A(puf_21_wire_8), .Y(outData[10]));
   BUFX2 puf_out_instance_21 ( .A(outData[10]), .Y(pufout[21]));
   INVX1 puf_22_instance_0 ( .A(puf_22_wire_1), .Y(puf_22_wire_0));
   MUX2X1 puf_22_instance_1 ( .A(puf_22_wire_0),  .B(outData[9]),  .S(sel), .Y(puf_22_wire_2));
   INVX1 puf_22_instance_2 ( .A(puf_22_wire_2), .Y(puf_22_wire_5));
   INVX1 puf_22_instance_3 ( .A(puf_22_wire_5), .Y(puf_22_wire_6));
   MUX2X1 puf_22_instance_4 ( .A(puf_22_wire_0),  .B(puf_22_wire_6),  .S(sel), .Y(puf_22_wire_7));
   INVX1 puf_22_instance_5 ( .A(puf_22_wire_7), .Y(puf_22_wire_8));
   INVX1 puf_22_instance_6 ( .A(puf_22_wire_8), .Y(outData[9]));
   BUFX2 puf_out_instance_22 ( .A(outData[9]), .Y(pufout[22]));
   INVX1 puf_23_instance_0 ( .A(puf_23_wire_1), .Y(puf_23_wire_0));
   MUX2X1 puf_23_instance_1 ( .A(puf_23_wire_0),  .B(outData[8]),  .S(sel), .Y(puf_23_wire_2));
   INVX1 puf_23_instance_2 ( .A(puf_23_wire_2), .Y(puf_23_wire_5));
   INVX1 puf_23_instance_3 ( .A(puf_23_wire_5), .Y(puf_23_wire_6));
   MUX2X1 puf_23_instance_4 ( .A(puf_23_wire_0),  .B(puf_23_wire_6),  .S(sel), .Y(puf_23_wire_7));
   INVX1 puf_23_instance_5 ( .A(puf_23_wire_7), .Y(puf_23_wire_8));
   INVX1 puf_23_instance_6 ( .A(puf_23_wire_8), .Y(outData[8]));
   BUFX2 puf_out_instance_23 ( .A(outData[8]), .Y(pufout[23]));
   INVX1 puf_24_instance_0 ( .A(puf_24_wire_1), .Y(puf_24_wire_0));
   MUX2X1 puf_24_instance_1 ( .A(puf_24_wire_0),  .B(outData[7]),  .S(sel), .Y(puf_24_wire_2));
   INVX1 puf_24_instance_2 ( .A(puf_24_wire_2), .Y(puf_24_wire_5));
   INVX1 puf_24_instance_3 ( .A(puf_24_wire_5), .Y(puf_24_wire_6));
   MUX2X1 puf_24_instance_4 ( .A(puf_24_wire_0),  .B(puf_24_wire_6),  .S(sel), .Y(puf_24_wire_7));
   INVX1 puf_24_instance_5 ( .A(puf_24_wire_7), .Y(puf_24_wire_8));
   INVX1 puf_24_instance_6 ( .A(puf_24_wire_8), .Y(outData[7]));
   BUFX2 puf_out_instance_24 ( .A(outData[7]), .Y(pufout[24]));
   INVX1 puf_25_instance_0 ( .A(puf_25_wire_1), .Y(puf_25_wire_0));
   MUX2X1 puf_25_instance_1 ( .A(puf_25_wire_0),  .B(outData[6]),  .S(sel), .Y(puf_25_wire_2));
   INVX1 puf_25_instance_2 ( .A(puf_25_wire_2), .Y(puf_25_wire_5));
   INVX1 puf_25_instance_3 ( .A(puf_25_wire_5), .Y(puf_25_wire_6));
   MUX2X1 puf_25_instance_4 ( .A(puf_25_wire_0),  .B(puf_25_wire_6),  .S(sel), .Y(puf_25_wire_7));
   INVX1 puf_25_instance_5 ( .A(puf_25_wire_7), .Y(puf_25_wire_8));
   INVX1 puf_25_instance_6 ( .A(puf_25_wire_8), .Y(outData[6]));
   BUFX2 puf_out_instance_25 ( .A(outData[6]), .Y(pufout[25]));
   INVX1 puf_26_instance_0 ( .A(puf_26_wire_1), .Y(puf_26_wire_0));
   MUX2X1 puf_26_instance_1 ( .A(puf_26_wire_0),  .B(outData[5]),  .S(sel), .Y(puf_26_wire_2));
   INVX1 puf_26_instance_2 ( .A(puf_26_wire_2), .Y(puf_26_wire_5));
   INVX1 puf_26_instance_3 ( .A(puf_26_wire_5), .Y(puf_26_wire_6));
   MUX2X1 puf_26_instance_4 ( .A(puf_26_wire_0),  .B(puf_26_wire_6),  .S(sel), .Y(puf_26_wire_7));
   INVX1 puf_26_instance_5 ( .A(puf_26_wire_7), .Y(puf_26_wire_8));
   INVX1 puf_26_instance_6 ( .A(puf_26_wire_8), .Y(outData[5]));
   BUFX2 puf_out_instance_26 ( .A(outData[5]), .Y(pufout[26]));
   INVX1 puf_27_instance_0 ( .A(puf_27_wire_1), .Y(puf_27_wire_0));
   MUX2X1 puf_27_instance_1 ( .A(puf_27_wire_0),  .B(outData[4]),  .S(sel), .Y(puf_27_wire_2));
   INVX1 puf_27_instance_2 ( .A(puf_27_wire_2), .Y(puf_27_wire_5));
   INVX1 puf_27_instance_3 ( .A(puf_27_wire_5), .Y(puf_27_wire_6));
   MUX2X1 puf_27_instance_4 ( .A(puf_27_wire_0),  .B(puf_27_wire_6),  .S(sel), .Y(puf_27_wire_7));
   INVX1 puf_27_instance_5 ( .A(puf_27_wire_7), .Y(puf_27_wire_8));
   INVX1 puf_27_instance_6 ( .A(puf_27_wire_8), .Y(outData[4]));
   BUFX2 puf_out_instance_27 ( .A(outData[4]), .Y(pufout[27]));
   INVX1 puf_28_instance_0 ( .A(puf_28_wire_1), .Y(puf_28_wire_0));
   MUX2X1 puf_28_instance_1 ( .A(puf_28_wire_0),  .B(outData[3]),  .S(sel), .Y(puf_28_wire_2));
   INVX1 puf_28_instance_2 ( .A(puf_28_wire_2), .Y(puf_28_wire_5));
   INVX1 puf_28_instance_3 ( .A(puf_28_wire_5), .Y(puf_28_wire_6));
   MUX2X1 puf_28_instance_4 ( .A(puf_28_wire_0),  .B(puf_28_wire_6),  .S(sel), .Y(puf_28_wire_7));
   INVX1 puf_28_instance_5 ( .A(puf_28_wire_7), .Y(puf_28_wire_8));
   INVX1 puf_28_instance_6 ( .A(puf_28_wire_8), .Y(outData[3]));
   BUFX2 puf_out_instance_28 ( .A(outData[3]), .Y(pufout[28]));
   INVX1 puf_29_instance_0 ( .A(puf_29_wire_1), .Y(puf_29_wire_0));
   MUX2X1 puf_29_instance_1 ( .A(puf_29_wire_0),  .B(outData[2]),  .S(sel), .Y(puf_29_wire_2));
   INVX1 puf_29_instance_2 ( .A(puf_29_wire_2), .Y(puf_29_wire_5));
   INVX1 puf_29_instance_3 ( .A(puf_29_wire_5), .Y(puf_29_wire_6));
   MUX2X1 puf_29_instance_4 ( .A(puf_29_wire_0),  .B(puf_29_wire_6),  .S(sel), .Y(puf_29_wire_7));
   INVX1 puf_29_instance_5 ( .A(puf_29_wire_7), .Y(puf_29_wire_8));
   INVX1 puf_29_instance_6 ( .A(puf_29_wire_8), .Y(outData[2]));
   BUFX2 puf_out_instance_29 ( .A(outData[2]), .Y(pufout[29]));
   INVX1 puf_30_instance_0 ( .A(puf_30_wire_1), .Y(puf_30_wire_0));
   MUX2X1 puf_30_instance_1 ( .A(puf_30_wire_0),  .B(outData[1]),  .S(sel), .Y(puf_30_wire_2));
   INVX1 puf_30_instance_2 ( .A(puf_30_wire_2), .Y(puf_30_wire_5));
   INVX1 puf_30_instance_3 ( .A(puf_30_wire_5), .Y(puf_30_wire_6));
   MUX2X1 puf_30_instance_4 ( .A(puf_30_wire_0),  .B(puf_30_wire_6),  .S(sel), .Y(puf_30_wire_7));
   INVX1 puf_30_instance_5 ( .A(puf_30_wire_7), .Y(puf_30_wire_8));
   INVX1 puf_30_instance_6 ( .A(puf_30_wire_8), .Y(outData[1]));
   BUFX2 puf_out_instance_30 ( .A(outData[1]), .Y(pufout[30]));
   INVX1 puf_31_instance_0 ( .A(puf_31_wire_1), .Y(puf_31_wire_0));
   MUX2X1 puf_31_instance_1 ( .A(puf_31_wire_0),  .B(outData[0]),  .S(sel), .Y(puf_31_wire_2));
   INVX1 puf_31_instance_2 ( .A(puf_31_wire_2), .Y(puf_31_wire_5));
   INVX1 puf_31_instance_3 ( .A(puf_31_wire_5), .Y(puf_31_wire_6));
   MUX2X1 puf_31_instance_4 ( .A(puf_31_wire_0),  .B(puf_31_wire_6),  .S(sel), .Y(puf_31_wire_7));
   INVX1 puf_31_instance_5 ( .A(puf_31_wire_7), .Y(puf_31_wire_8));
   INVX1 puf_31_instance_6 ( .A(puf_31_wire_8), .Y(outData[0]));
   BUFX2 puf_out_instance_31 ( .A(outData[0]), .Y(pufout[31]));
   INVX1 puf_32_instance_0 ( .A(puf_32_wire_1), .Y(puf_32_wire_0));
   MUX2X1 puf_32_instance_1 ( .A(puf_32_wire_0),  .B(my_FIR_filter_firBlock_left_Y_in_0_),  .S(sel), .Y(puf_32_wire_2));
   INVX1 puf_32_instance_2 ( .A(puf_32_wire_2), .Y(puf_32_wire_5));
   INVX1 puf_32_instance_3 ( .A(puf_32_wire_5), .Y(puf_32_wire_6));
   MUX2X1 puf_32_instance_4 ( .A(puf_32_wire_0),  .B(puf_32_wire_6),  .S(sel), .Y(puf_32_wire_7));
   INVX1 puf_32_instance_5 ( .A(puf_32_wire_7), .Y(puf_32_wire_8));
   INVX1 puf_32_instance_6 ( .A(puf_32_wire_8), .Y(my_FIR_filter_firBlock_left_Y_in_0_));
   BUFX2 puf_out_instance_32 ( .A(my_FIR_filter_firBlock_left_Y_in_0_), .Y(pufout[32]));
   INVX1 puf_33_instance_0 ( .A(puf_33_wire_1), .Y(puf_33_wire_0));
   MUX2X1 puf_33_instance_1 ( .A(puf_33_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[0]),  .S(sel), .Y(puf_33_wire_2));
   INVX1 puf_33_instance_2 ( .A(puf_33_wire_2), .Y(puf_33_wire_5));
   INVX1 puf_33_instance_3 ( .A(puf_33_wire_5), .Y(puf_33_wire_6));
   MUX2X1 puf_33_instance_4 ( .A(puf_33_wire_0),  .B(puf_33_wire_6),  .S(sel), .Y(puf_33_wire_7));
   INVX1 puf_33_instance_5 ( .A(puf_33_wire_7), .Y(puf_33_wire_8));
   INVX1 puf_33_instance_6 ( .A(puf_33_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[0]));
   BUFX2 puf_out_instance_33 ( .A(my_FIR_filter_firBlock_left_firStep[0]), .Y(pufout[33]));
   INVX1 puf_34_instance_0 ( .A(puf_34_wire_1), .Y(puf_34_wire_0));
   MUX2X1 puf_34_instance_1 ( .A(puf_34_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[1]),  .S(sel), .Y(puf_34_wire_2));
   INVX1 puf_34_instance_2 ( .A(puf_34_wire_2), .Y(puf_34_wire_5));
   INVX1 puf_34_instance_3 ( .A(puf_34_wire_5), .Y(puf_34_wire_6));
   MUX2X1 puf_34_instance_4 ( .A(puf_34_wire_0),  .B(puf_34_wire_6),  .S(sel), .Y(puf_34_wire_7));
   INVX1 puf_34_instance_5 ( .A(puf_34_wire_7), .Y(puf_34_wire_8));
   INVX1 puf_34_instance_6 ( .A(puf_34_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[1]));
   BUFX2 puf_out_instance_34 ( .A(my_FIR_filter_firBlock_left_firStep[1]), .Y(pufout[34]));
   INVX1 puf_35_instance_0 ( .A(puf_35_wire_1), .Y(puf_35_wire_0));
   MUX2X1 puf_35_instance_1 ( .A(puf_35_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[2]),  .S(sel), .Y(puf_35_wire_2));
   INVX1 puf_35_instance_2 ( .A(puf_35_wire_2), .Y(puf_35_wire_5));
   INVX1 puf_35_instance_3 ( .A(puf_35_wire_5), .Y(puf_35_wire_6));
   MUX2X1 puf_35_instance_4 ( .A(puf_35_wire_0),  .B(puf_35_wire_6),  .S(sel), .Y(puf_35_wire_7));
   INVX1 puf_35_instance_5 ( .A(puf_35_wire_7), .Y(puf_35_wire_8));
   INVX1 puf_35_instance_6 ( .A(puf_35_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[2]));
   BUFX2 puf_out_instance_35 ( .A(my_FIR_filter_firBlock_left_firStep[2]), .Y(pufout[35]));
   INVX1 puf_36_instance_0 ( .A(puf_36_wire_1), .Y(puf_36_wire_0));
   MUX2X1 puf_36_instance_1 ( .A(puf_36_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[3]),  .S(sel), .Y(puf_36_wire_2));
   INVX1 puf_36_instance_2 ( .A(puf_36_wire_2), .Y(puf_36_wire_5));
   INVX1 puf_36_instance_3 ( .A(puf_36_wire_5), .Y(puf_36_wire_6));
   MUX2X1 puf_36_instance_4 ( .A(puf_36_wire_0),  .B(puf_36_wire_6),  .S(sel), .Y(puf_36_wire_7));
   INVX1 puf_36_instance_5 ( .A(puf_36_wire_7), .Y(puf_36_wire_8));
   INVX1 puf_36_instance_6 ( .A(puf_36_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[3]));
   BUFX2 puf_out_instance_36 ( .A(my_FIR_filter_firBlock_left_firStep[3]), .Y(pufout[36]));
   INVX1 puf_37_instance_0 ( .A(puf_37_wire_1), .Y(puf_37_wire_0));
   MUX2X1 puf_37_instance_1 ( .A(puf_37_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[4]),  .S(sel), .Y(puf_37_wire_2));
   INVX1 puf_37_instance_2 ( .A(puf_37_wire_2), .Y(puf_37_wire_5));
   INVX1 puf_37_instance_3 ( .A(puf_37_wire_5), .Y(puf_37_wire_6));
   MUX2X1 puf_37_instance_4 ( .A(puf_37_wire_0),  .B(puf_37_wire_6),  .S(sel), .Y(puf_37_wire_7));
   INVX1 puf_37_instance_5 ( .A(puf_37_wire_7), .Y(puf_37_wire_8));
   INVX1 puf_37_instance_6 ( .A(puf_37_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[4]));
   BUFX2 puf_out_instance_37 ( .A(my_FIR_filter_firBlock_left_firStep[4]), .Y(pufout[37]));
   INVX1 puf_38_instance_0 ( .A(puf_38_wire_1), .Y(puf_38_wire_0));
   MUX2X1 puf_38_instance_1 ( .A(puf_38_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[5]),  .S(sel), .Y(puf_38_wire_2));
   INVX1 puf_38_instance_2 ( .A(puf_38_wire_2), .Y(puf_38_wire_5));
   INVX1 puf_38_instance_3 ( .A(puf_38_wire_5), .Y(puf_38_wire_6));
   MUX2X1 puf_38_instance_4 ( .A(puf_38_wire_0),  .B(puf_38_wire_6),  .S(sel), .Y(puf_38_wire_7));
   INVX1 puf_38_instance_5 ( .A(puf_38_wire_7), .Y(puf_38_wire_8));
   INVX1 puf_38_instance_6 ( .A(puf_38_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[5]));
   BUFX2 puf_out_instance_38 ( .A(my_FIR_filter_firBlock_left_firStep[5]), .Y(pufout[38]));
   INVX1 puf_39_instance_0 ( .A(puf_39_wire_1), .Y(puf_39_wire_0));
   MUX2X1 puf_39_instance_1 ( .A(puf_39_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[6]),  .S(sel), .Y(puf_39_wire_2));
   INVX1 puf_39_instance_2 ( .A(puf_39_wire_2), .Y(puf_39_wire_5));
   INVX1 puf_39_instance_3 ( .A(puf_39_wire_5), .Y(puf_39_wire_6));
   MUX2X1 puf_39_instance_4 ( .A(puf_39_wire_0),  .B(puf_39_wire_6),  .S(sel), .Y(puf_39_wire_7));
   INVX1 puf_39_instance_5 ( .A(puf_39_wire_7), .Y(puf_39_wire_8));
   INVX1 puf_39_instance_6 ( .A(puf_39_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[6]));
   BUFX2 puf_out_instance_39 ( .A(my_FIR_filter_firBlock_left_firStep[6]), .Y(pufout[39]));
   INVX1 puf_40_instance_0 ( .A(puf_40_wire_1), .Y(puf_40_wire_0));
   MUX2X1 puf_40_instance_1 ( .A(puf_40_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[7]),  .S(sel), .Y(puf_40_wire_2));
   INVX1 puf_40_instance_2 ( .A(puf_40_wire_2), .Y(puf_40_wire_5));
   INVX1 puf_40_instance_3 ( .A(puf_40_wire_5), .Y(puf_40_wire_6));
   MUX2X1 puf_40_instance_4 ( .A(puf_40_wire_0),  .B(puf_40_wire_6),  .S(sel), .Y(puf_40_wire_7));
   INVX1 puf_40_instance_5 ( .A(puf_40_wire_7), .Y(puf_40_wire_8));
   INVX1 puf_40_instance_6 ( .A(puf_40_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[7]));
   BUFX2 puf_out_instance_40 ( .A(my_FIR_filter_firBlock_left_firStep[7]), .Y(pufout[40]));
   INVX1 puf_41_instance_0 ( .A(puf_41_wire_1), .Y(puf_41_wire_0));
   MUX2X1 puf_41_instance_1 ( .A(puf_41_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[8]),  .S(sel), .Y(puf_41_wire_2));
   INVX1 puf_41_instance_2 ( .A(puf_41_wire_2), .Y(puf_41_wire_5));
   INVX1 puf_41_instance_3 ( .A(puf_41_wire_5), .Y(puf_41_wire_6));
   MUX2X1 puf_41_instance_4 ( .A(puf_41_wire_0),  .B(puf_41_wire_6),  .S(sel), .Y(puf_41_wire_7));
   INVX1 puf_41_instance_5 ( .A(puf_41_wire_7), .Y(puf_41_wire_8));
   INVX1 puf_41_instance_6 ( .A(puf_41_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[8]));
   BUFX2 puf_out_instance_41 ( .A(my_FIR_filter_firBlock_left_firStep[8]), .Y(pufout[41]));
   INVX1 puf_42_instance_0 ( .A(puf_42_wire_1), .Y(puf_42_wire_0));
   MUX2X1 puf_42_instance_1 ( .A(puf_42_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[9]),  .S(sel), .Y(puf_42_wire_2));
   INVX1 puf_42_instance_2 ( .A(puf_42_wire_2), .Y(puf_42_wire_5));
   INVX1 puf_42_instance_3 ( .A(puf_42_wire_5), .Y(puf_42_wire_6));
   MUX2X1 puf_42_instance_4 ( .A(puf_42_wire_0),  .B(puf_42_wire_6),  .S(sel), .Y(puf_42_wire_7));
   INVX1 puf_42_instance_5 ( .A(puf_42_wire_7), .Y(puf_42_wire_8));
   INVX1 puf_42_instance_6 ( .A(puf_42_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[9]));
   BUFX2 puf_out_instance_42 ( .A(my_FIR_filter_firBlock_left_firStep[9]), .Y(pufout[42]));
   INVX1 puf_43_instance_0 ( .A(puf_43_wire_1), .Y(puf_43_wire_0));
   MUX2X1 puf_43_instance_1 ( .A(puf_43_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[10]),  .S(sel), .Y(puf_43_wire_2));
   INVX1 puf_43_instance_2 ( .A(puf_43_wire_2), .Y(puf_43_wire_5));
   INVX1 puf_43_instance_3 ( .A(puf_43_wire_5), .Y(puf_43_wire_6));
   MUX2X1 puf_43_instance_4 ( .A(puf_43_wire_0),  .B(puf_43_wire_6),  .S(sel), .Y(puf_43_wire_7));
   INVX1 puf_43_instance_5 ( .A(puf_43_wire_7), .Y(puf_43_wire_8));
   INVX1 puf_43_instance_6 ( .A(puf_43_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[10]));
   BUFX2 puf_out_instance_43 ( .A(my_FIR_filter_firBlock_left_firStep[10]), .Y(pufout[43]));
   INVX1 puf_44_instance_0 ( .A(puf_44_wire_1), .Y(puf_44_wire_0));
   MUX2X1 puf_44_instance_1 ( .A(puf_44_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[11]),  .S(sel), .Y(puf_44_wire_2));
   INVX1 puf_44_instance_2 ( .A(puf_44_wire_2), .Y(puf_44_wire_5));
   INVX1 puf_44_instance_3 ( .A(puf_44_wire_5), .Y(puf_44_wire_6));
   MUX2X1 puf_44_instance_4 ( .A(puf_44_wire_0),  .B(puf_44_wire_6),  .S(sel), .Y(puf_44_wire_7));
   INVX1 puf_44_instance_5 ( .A(puf_44_wire_7), .Y(puf_44_wire_8));
   INVX1 puf_44_instance_6 ( .A(puf_44_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[11]));
   BUFX2 puf_out_instance_44 ( .A(my_FIR_filter_firBlock_left_firStep[11]), .Y(pufout[44]));
   INVX1 puf_45_instance_0 ( .A(puf_45_wire_1), .Y(puf_45_wire_0));
   MUX2X1 puf_45_instance_1 ( .A(puf_45_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[12]),  .S(sel), .Y(puf_45_wire_2));
   INVX1 puf_45_instance_2 ( .A(puf_45_wire_2), .Y(puf_45_wire_5));
   INVX1 puf_45_instance_3 ( .A(puf_45_wire_5), .Y(puf_45_wire_6));
   MUX2X1 puf_45_instance_4 ( .A(puf_45_wire_0),  .B(puf_45_wire_6),  .S(sel), .Y(puf_45_wire_7));
   INVX1 puf_45_instance_5 ( .A(puf_45_wire_7), .Y(puf_45_wire_8));
   INVX1 puf_45_instance_6 ( .A(puf_45_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[12]));
   BUFX2 puf_out_instance_45 ( .A(my_FIR_filter_firBlock_left_firStep[12]), .Y(pufout[45]));
   INVX1 puf_46_instance_0 ( .A(puf_46_wire_1), .Y(puf_46_wire_0));
   MUX2X1 puf_46_instance_1 ( .A(puf_46_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[13]),  .S(sel), .Y(puf_46_wire_2));
   INVX1 puf_46_instance_2 ( .A(puf_46_wire_2), .Y(puf_46_wire_5));
   INVX1 puf_46_instance_3 ( .A(puf_46_wire_5), .Y(puf_46_wire_6));
   MUX2X1 puf_46_instance_4 ( .A(puf_46_wire_0),  .B(puf_46_wire_6),  .S(sel), .Y(puf_46_wire_7));
   INVX1 puf_46_instance_5 ( .A(puf_46_wire_7), .Y(puf_46_wire_8));
   INVX1 puf_46_instance_6 ( .A(puf_46_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[13]));
   BUFX2 puf_out_instance_46 ( .A(my_FIR_filter_firBlock_left_firStep[13]), .Y(pufout[46]));
   INVX1 puf_47_instance_0 ( .A(puf_47_wire_1), .Y(puf_47_wire_0));
   MUX2X1 puf_47_instance_1 ( .A(puf_47_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[14]),  .S(sel), .Y(puf_47_wire_2));
   INVX1 puf_47_instance_2 ( .A(puf_47_wire_2), .Y(puf_47_wire_5));
   INVX1 puf_47_instance_3 ( .A(puf_47_wire_5), .Y(puf_47_wire_6));
   MUX2X1 puf_47_instance_4 ( .A(puf_47_wire_0),  .B(puf_47_wire_6),  .S(sel), .Y(puf_47_wire_7));
   INVX1 puf_47_instance_5 ( .A(puf_47_wire_7), .Y(puf_47_wire_8));
   INVX1 puf_47_instance_6 ( .A(puf_47_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[14]));
   BUFX2 puf_out_instance_47 ( .A(my_FIR_filter_firBlock_left_firStep[14]), .Y(pufout[47]));
   INVX1 puf_48_instance_0 ( .A(puf_48_wire_1), .Y(puf_48_wire_0));
   MUX2X1 puf_48_instance_1 ( .A(puf_48_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[15]),  .S(sel), .Y(puf_48_wire_2));
   INVX1 puf_48_instance_2 ( .A(puf_48_wire_2), .Y(puf_48_wire_5));
   INVX1 puf_48_instance_3 ( .A(puf_48_wire_5), .Y(puf_48_wire_6));
   MUX2X1 puf_48_instance_4 ( .A(puf_48_wire_0),  .B(puf_48_wire_6),  .S(sel), .Y(puf_48_wire_7));
   INVX1 puf_48_instance_5 ( .A(puf_48_wire_7), .Y(puf_48_wire_8));
   INVX1 puf_48_instance_6 ( .A(puf_48_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[15]));
   BUFX2 puf_out_instance_48 ( .A(my_FIR_filter_firBlock_left_firStep[15]), .Y(pufout[48]));
   INVX1 puf_49_instance_0 ( .A(puf_49_wire_1), .Y(puf_49_wire_0));
   MUX2X1 puf_49_instance_1 ( .A(puf_49_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[16]),  .S(sel), .Y(puf_49_wire_2));
   INVX1 puf_49_instance_2 ( .A(puf_49_wire_2), .Y(puf_49_wire_5));
   INVX1 puf_49_instance_3 ( .A(puf_49_wire_5), .Y(puf_49_wire_6));
   MUX2X1 puf_49_instance_4 ( .A(puf_49_wire_0),  .B(puf_49_wire_6),  .S(sel), .Y(puf_49_wire_7));
   INVX1 puf_49_instance_5 ( .A(puf_49_wire_7), .Y(puf_49_wire_8));
   INVX1 puf_49_instance_6 ( .A(puf_49_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[16]));
   BUFX2 puf_out_instance_49 ( .A(my_FIR_filter_firBlock_left_firStep[16]), .Y(pufout[49]));
   INVX1 puf_50_instance_0 ( .A(puf_50_wire_1), .Y(puf_50_wire_0));
   MUX2X1 puf_50_instance_1 ( .A(puf_50_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[17]),  .S(sel), .Y(puf_50_wire_2));
   INVX1 puf_50_instance_2 ( .A(puf_50_wire_2), .Y(puf_50_wire_5));
   INVX1 puf_50_instance_3 ( .A(puf_50_wire_5), .Y(puf_50_wire_6));
   MUX2X1 puf_50_instance_4 ( .A(puf_50_wire_0),  .B(puf_50_wire_6),  .S(sel), .Y(puf_50_wire_7));
   INVX1 puf_50_instance_5 ( .A(puf_50_wire_7), .Y(puf_50_wire_8));
   INVX1 puf_50_instance_6 ( .A(puf_50_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[17]));
   BUFX2 puf_out_instance_50 ( .A(my_FIR_filter_firBlock_left_firStep[17]), .Y(pufout[50]));
   INVX1 puf_51_instance_0 ( .A(puf_51_wire_1), .Y(puf_51_wire_0));
   MUX2X1 puf_51_instance_1 ( .A(puf_51_wire_0),  .B(my_FIR_filter_firBlock_left_firStep[18]),  .S(sel), .Y(puf_51_wire_2));
   INVX1 puf_51_instance_2 ( .A(puf_51_wire_2), .Y(puf_51_wire_5));
   INVX1 puf_51_instance_3 ( .A(puf_51_wire_5), .Y(puf_51_wire_6));
   MUX2X1 puf_51_instance_4 ( .A(puf_51_wire_0),  .B(puf_51_wire_6),  .S(sel), .Y(puf_51_wire_7));
   INVX1 puf_51_instance_5 ( .A(puf_51_wire_7), .Y(puf_51_wire_8));
   INVX1 puf_51_instance_6 ( .A(puf_51_wire_8), .Y(my_FIR_filter_firBlock_left_firStep[18]));
   BUFX2 puf_out_instance_51 ( .A(my_FIR_filter_firBlock_left_firStep[18]), .Y(pufout[51]));
   INVX1 puf_52_instance_0 ( .A(puf_52_wire_1), .Y(puf_52_wire_0));
   MUX2X1 puf_52_instance_1 ( .A(puf_52_wire_0),  .B(n67),  .S(sel), .Y(puf_52_wire_2));
   INVX1 puf_52_instance_2 ( .A(puf_52_wire_2), .Y(puf_52_wire_5));
   INVX1 puf_52_instance_3 ( .A(puf_52_wire_5), .Y(puf_52_wire_6));
   MUX2X1 puf_52_instance_4 ( .A(puf_52_wire_0),  .B(puf_52_wire_6),  .S(sel), .Y(puf_52_wire_7));
   INVX1 puf_52_instance_5 ( .A(puf_52_wire_7), .Y(puf_52_wire_8));
   INVX1 puf_52_instance_6 ( .A(puf_52_wire_8), .Y(n67));
   BUFX2 puf_out_instance_52 ( .A(n67), .Y(pufout[52]));
   INVX1 puf_53_instance_0 ( .A(puf_53_wire_1), .Y(puf_53_wire_0));
   MUX2X1 puf_53_instance_1 ( .A(puf_53_wire_0),  .B(n68),  .S(sel), .Y(puf_53_wire_2));
   INVX1 puf_53_instance_2 ( .A(puf_53_wire_2), .Y(puf_53_wire_5));
   INVX1 puf_53_instance_3 ( .A(puf_53_wire_5), .Y(puf_53_wire_6));
   MUX2X1 puf_53_instance_4 ( .A(puf_53_wire_0),  .B(puf_53_wire_6),  .S(sel), .Y(puf_53_wire_7));
   INVX1 puf_53_instance_5 ( .A(puf_53_wire_7), .Y(puf_53_wire_8));
   INVX1 puf_53_instance_6 ( .A(puf_53_wire_8), .Y(n68));
   BUFX2 puf_out_instance_53 ( .A(n68), .Y(pufout[53]));
   INVX1 puf_54_instance_0 ( .A(puf_54_wire_1), .Y(puf_54_wire_0));
   MUX2X1 puf_54_instance_1 ( .A(puf_54_wire_0),  .B(n69),  .S(sel), .Y(puf_54_wire_2));
   INVX1 puf_54_instance_2 ( .A(puf_54_wire_2), .Y(puf_54_wire_5));
   INVX1 puf_54_instance_3 ( .A(puf_54_wire_5), .Y(puf_54_wire_6));
   MUX2X1 puf_54_instance_4 ( .A(puf_54_wire_0),  .B(puf_54_wire_6),  .S(sel), .Y(puf_54_wire_7));
   INVX1 puf_54_instance_5 ( .A(puf_54_wire_7), .Y(puf_54_wire_8));
   INVX1 puf_54_instance_6 ( .A(puf_54_wire_8), .Y(n69));
   BUFX2 puf_out_instance_54 ( .A(n69), .Y(pufout[54]));
   INVX1 puf_55_instance_0 ( .A(puf_55_wire_1), .Y(puf_55_wire_0));
   MUX2X1 puf_55_instance_1 ( .A(puf_55_wire_0),  .B(n70),  .S(sel), .Y(puf_55_wire_2));
   INVX1 puf_55_instance_2 ( .A(puf_55_wire_2), .Y(puf_55_wire_5));
   INVX1 puf_55_instance_3 ( .A(puf_55_wire_5), .Y(puf_55_wire_6));
   MUX2X1 puf_55_instance_4 ( .A(puf_55_wire_0),  .B(puf_55_wire_6),  .S(sel), .Y(puf_55_wire_7));
   INVX1 puf_55_instance_5 ( .A(puf_55_wire_7), .Y(puf_55_wire_8));
   INVX1 puf_55_instance_6 ( .A(puf_55_wire_8), .Y(n70));
   BUFX2 puf_out_instance_55 ( .A(n70), .Y(pufout[55]));
   INVX1 puf_56_instance_0 ( .A(puf_56_wire_1), .Y(puf_56_wire_0));
   MUX2X1 puf_56_instance_1 ( .A(puf_56_wire_0),  .B(n71),  .S(sel), .Y(puf_56_wire_2));
   INVX1 puf_56_instance_2 ( .A(puf_56_wire_2), .Y(puf_56_wire_5));
   INVX1 puf_56_instance_3 ( .A(puf_56_wire_5), .Y(puf_56_wire_6));
   MUX2X1 puf_56_instance_4 ( .A(puf_56_wire_0),  .B(puf_56_wire_6),  .S(sel), .Y(puf_56_wire_7));
   INVX1 puf_56_instance_5 ( .A(puf_56_wire_7), .Y(puf_56_wire_8));
   INVX1 puf_56_instance_6 ( .A(puf_56_wire_8), .Y(n71));
   BUFX2 puf_out_instance_56 ( .A(n71), .Y(pufout[56]));
   INVX1 puf_57_instance_0 ( .A(puf_57_wire_1), .Y(puf_57_wire_0));
   MUX2X1 puf_57_instance_1 ( .A(puf_57_wire_0),  .B(n72),  .S(sel), .Y(puf_57_wire_2));
   INVX1 puf_57_instance_2 ( .A(puf_57_wire_2), .Y(puf_57_wire_5));
   INVX1 puf_57_instance_3 ( .A(puf_57_wire_5), .Y(puf_57_wire_6));
   MUX2X1 puf_57_instance_4 ( .A(puf_57_wire_0),  .B(puf_57_wire_6),  .S(sel), .Y(puf_57_wire_7));
   INVX1 puf_57_instance_5 ( .A(puf_57_wire_7), .Y(puf_57_wire_8));
   INVX1 puf_57_instance_6 ( .A(puf_57_wire_8), .Y(n72));
   BUFX2 puf_out_instance_57 ( .A(n72), .Y(pufout[57]));
   INVX1 puf_58_instance_0 ( .A(puf_58_wire_1), .Y(puf_58_wire_0));
   MUX2X1 puf_58_instance_1 ( .A(puf_58_wire_0),  .B(n73),  .S(sel), .Y(puf_58_wire_2));
   INVX1 puf_58_instance_2 ( .A(puf_58_wire_2), .Y(puf_58_wire_5));
   INVX1 puf_58_instance_3 ( .A(puf_58_wire_5), .Y(puf_58_wire_6));
   MUX2X1 puf_58_instance_4 ( .A(puf_58_wire_0),  .B(puf_58_wire_6),  .S(sel), .Y(puf_58_wire_7));
   INVX1 puf_58_instance_5 ( .A(puf_58_wire_7), .Y(puf_58_wire_8));
   INVX1 puf_58_instance_6 ( .A(puf_58_wire_8), .Y(n73));
   BUFX2 puf_out_instance_58 ( .A(n73), .Y(pufout[58]));
   INVX1 puf_59_instance_0 ( .A(puf_59_wire_1), .Y(puf_59_wire_0));
   MUX2X1 puf_59_instance_1 ( .A(puf_59_wire_0),  .B(n74),  .S(sel), .Y(puf_59_wire_2));
   INVX1 puf_59_instance_2 ( .A(puf_59_wire_2), .Y(puf_59_wire_5));
   INVX1 puf_59_instance_3 ( .A(puf_59_wire_5), .Y(puf_59_wire_6));
   MUX2X1 puf_59_instance_4 ( .A(puf_59_wire_0),  .B(puf_59_wire_6),  .S(sel), .Y(puf_59_wire_7));
   INVX1 puf_59_instance_5 ( .A(puf_59_wire_7), .Y(puf_59_wire_8));
   INVX1 puf_59_instance_6 ( .A(puf_59_wire_8), .Y(n74));
   BUFX2 puf_out_instance_59 ( .A(n74), .Y(pufout[59]));
   INVX1 puf_60_instance_0 ( .A(puf_60_wire_1), .Y(puf_60_wire_0));
   MUX2X1 puf_60_instance_1 ( .A(puf_60_wire_0),  .B(n75),  .S(sel), .Y(puf_60_wire_2));
   INVX1 puf_60_instance_2 ( .A(puf_60_wire_2), .Y(puf_60_wire_5));
   INVX1 puf_60_instance_3 ( .A(puf_60_wire_5), .Y(puf_60_wire_6));
   MUX2X1 puf_60_instance_4 ( .A(puf_60_wire_0),  .B(puf_60_wire_6),  .S(sel), .Y(puf_60_wire_7));
   INVX1 puf_60_instance_5 ( .A(puf_60_wire_7), .Y(puf_60_wire_8));
   INVX1 puf_60_instance_6 ( .A(puf_60_wire_8), .Y(n75));
   BUFX2 puf_out_instance_60 ( .A(n75), .Y(pufout[60]));
   INVX1 puf_61_instance_0 ( .A(puf_61_wire_1), .Y(puf_61_wire_0));
   MUX2X1 puf_61_instance_1 ( .A(puf_61_wire_0),  .B(n76),  .S(sel), .Y(puf_61_wire_2));
   INVX1 puf_61_instance_2 ( .A(puf_61_wire_2), .Y(puf_61_wire_5));
   INVX1 puf_61_instance_3 ( .A(puf_61_wire_5), .Y(puf_61_wire_6));
   MUX2X1 puf_61_instance_4 ( .A(puf_61_wire_0),  .B(puf_61_wire_6),  .S(sel), .Y(puf_61_wire_7));
   INVX1 puf_61_instance_5 ( .A(puf_61_wire_7), .Y(puf_61_wire_8));
   INVX1 puf_61_instance_6 ( .A(puf_61_wire_8), .Y(n76));
   BUFX2 puf_out_instance_61 ( .A(n76), .Y(pufout[61]));
   INVX1 puf_62_instance_0 ( .A(puf_62_wire_1), .Y(puf_62_wire_0));
   MUX2X1 puf_62_instance_1 ( .A(puf_62_wire_0),  .B(n77),  .S(sel), .Y(puf_62_wire_2));
   INVX1 puf_62_instance_2 ( .A(puf_62_wire_2), .Y(puf_62_wire_5));
   INVX1 puf_62_instance_3 ( .A(puf_62_wire_5), .Y(puf_62_wire_6));
   MUX2X1 puf_62_instance_4 ( .A(puf_62_wire_0),  .B(puf_62_wire_6),  .S(sel), .Y(puf_62_wire_7));
   INVX1 puf_62_instance_5 ( .A(puf_62_wire_7), .Y(puf_62_wire_8));
   INVX1 puf_62_instance_6 ( .A(puf_62_wire_8), .Y(n77));
   BUFX2 puf_out_instance_62 ( .A(n77), .Y(pufout[62]));
   INVX1 puf_63_instance_0 ( .A(puf_63_wire_1), .Y(puf_63_wire_0));
   MUX2X1 puf_63_instance_1 ( .A(puf_63_wire_0),  .B(n78),  .S(sel), .Y(puf_63_wire_2));
   INVX1 puf_63_instance_2 ( .A(puf_63_wire_2), .Y(puf_63_wire_5));
   INVX1 puf_63_instance_3 ( .A(puf_63_wire_5), .Y(puf_63_wire_6));
   MUX2X1 puf_63_instance_4 ( .A(puf_63_wire_0),  .B(puf_63_wire_6),  .S(sel), .Y(puf_63_wire_7));
   INVX1 puf_63_instance_5 ( .A(puf_63_wire_7), .Y(puf_63_wire_8));
   INVX1 puf_63_instance_6 ( .A(puf_63_wire_8), .Y(n78));
   BUFX2 puf_out_instance_63 ( .A(n78), .Y(pufout[63]));
   INVX1 puf_64_instance_0 ( .A(puf_64_wire_1), .Y(puf_64_wire_0));
   MUX2X1 puf_64_instance_1 ( .A(puf_64_wire_0),  .B(n79),  .S(sel), .Y(puf_64_wire_2));
   INVX1 puf_64_instance_2 ( .A(puf_64_wire_2), .Y(puf_64_wire_5));
   INVX1 puf_64_instance_3 ( .A(puf_64_wire_5), .Y(puf_64_wire_6));
   MUX2X1 puf_64_instance_4 ( .A(puf_64_wire_0),  .B(puf_64_wire_6),  .S(sel), .Y(puf_64_wire_7));
   INVX1 puf_64_instance_5 ( .A(puf_64_wire_7), .Y(puf_64_wire_8));
   INVX1 puf_64_instance_6 ( .A(puf_64_wire_8), .Y(n79));
   BUFX2 puf_out_instance_64 ( .A(n79), .Y(pufout[64]));
   INVX1 puf_65_instance_0 ( .A(puf_65_wire_1), .Y(puf_65_wire_0));
   MUX2X1 puf_65_instance_1 ( .A(puf_65_wire_0),  .B(n80),  .S(sel), .Y(puf_65_wire_2));
   INVX1 puf_65_instance_2 ( .A(puf_65_wire_2), .Y(puf_65_wire_5));
   INVX1 puf_65_instance_3 ( .A(puf_65_wire_5), .Y(puf_65_wire_6));
   MUX2X1 puf_65_instance_4 ( .A(puf_65_wire_0),  .B(puf_65_wire_6),  .S(sel), .Y(puf_65_wire_7));
   INVX1 puf_65_instance_5 ( .A(puf_65_wire_7), .Y(puf_65_wire_8));
   INVX1 puf_65_instance_6 ( .A(puf_65_wire_8), .Y(n80));
   BUFX2 puf_out_instance_65 ( .A(n80), .Y(pufout[65]));
   INVX1 puf_66_instance_0 ( .A(puf_66_wire_1), .Y(puf_66_wire_0));
   MUX2X1 puf_66_instance_1 ( .A(puf_66_wire_0),  .B(n81),  .S(sel), .Y(puf_66_wire_2));
   INVX1 puf_66_instance_2 ( .A(puf_66_wire_2), .Y(puf_66_wire_5));
   INVX1 puf_66_instance_3 ( .A(puf_66_wire_5), .Y(puf_66_wire_6));
   MUX2X1 puf_66_instance_4 ( .A(puf_66_wire_0),  .B(puf_66_wire_6),  .S(sel), .Y(puf_66_wire_7));
   INVX1 puf_66_instance_5 ( .A(puf_66_wire_7), .Y(puf_66_wire_8));
   INVX1 puf_66_instance_6 ( .A(puf_66_wire_8), .Y(n81));
   BUFX2 puf_out_instance_66 ( .A(n81), .Y(pufout[66]));
   INVX1 puf_67_instance_0 ( .A(puf_67_wire_1), .Y(puf_67_wire_0));
   MUX2X1 puf_67_instance_1 ( .A(puf_67_wire_0),  .B(n82),  .S(sel), .Y(puf_67_wire_2));
   INVX1 puf_67_instance_2 ( .A(puf_67_wire_2), .Y(puf_67_wire_5));
   INVX1 puf_67_instance_3 ( .A(puf_67_wire_5), .Y(puf_67_wire_6));
   MUX2X1 puf_67_instance_4 ( .A(puf_67_wire_0),  .B(puf_67_wire_6),  .S(sel), .Y(puf_67_wire_7));
   INVX1 puf_67_instance_5 ( .A(puf_67_wire_7), .Y(puf_67_wire_8));
   INVX1 puf_67_instance_6 ( .A(puf_67_wire_8), .Y(n82));
   BUFX2 puf_out_instance_67 ( .A(n82), .Y(pufout[67]));
   INVX1 puf_68_instance_0 ( .A(puf_68_wire_1), .Y(puf_68_wire_0));
   MUX2X1 puf_68_instance_1 ( .A(puf_68_wire_0),  .B(n83),  .S(sel), .Y(puf_68_wire_2));
   INVX1 puf_68_instance_2 ( .A(puf_68_wire_2), .Y(puf_68_wire_5));
   INVX1 puf_68_instance_3 ( .A(puf_68_wire_5), .Y(puf_68_wire_6));
   MUX2X1 puf_68_instance_4 ( .A(puf_68_wire_0),  .B(puf_68_wire_6),  .S(sel), .Y(puf_68_wire_7));
   INVX1 puf_68_instance_5 ( .A(puf_68_wire_7), .Y(puf_68_wire_8));
   INVX1 puf_68_instance_6 ( .A(puf_68_wire_8), .Y(n83));
   BUFX2 puf_out_instance_68 ( .A(n83), .Y(pufout[68]));
   INVX1 puf_69_instance_0 ( .A(puf_69_wire_1), .Y(puf_69_wire_0));
   MUX2X1 puf_69_instance_1 ( .A(puf_69_wire_0),  .B(n84),  .S(sel), .Y(puf_69_wire_2));
   INVX1 puf_69_instance_2 ( .A(puf_69_wire_2), .Y(puf_69_wire_5));
   INVX1 puf_69_instance_3 ( .A(puf_69_wire_5), .Y(puf_69_wire_6));
   MUX2X1 puf_69_instance_4 ( .A(puf_69_wire_0),  .B(puf_69_wire_6),  .S(sel), .Y(puf_69_wire_7));
   INVX1 puf_69_instance_5 ( .A(puf_69_wire_7), .Y(puf_69_wire_8));
   INVX1 puf_69_instance_6 ( .A(puf_69_wire_8), .Y(n84));
   BUFX2 puf_out_instance_69 ( .A(n84), .Y(pufout[69]));
   INVX1 puf_70_instance_0 ( .A(puf_70_wire_1), .Y(puf_70_wire_0));
   MUX2X1 puf_70_instance_1 ( .A(puf_70_wire_0),  .B(n85),  .S(sel), .Y(puf_70_wire_2));
   INVX1 puf_70_instance_2 ( .A(puf_70_wire_2), .Y(puf_70_wire_5));
   INVX1 puf_70_instance_3 ( .A(puf_70_wire_5), .Y(puf_70_wire_6));
   MUX2X1 puf_70_instance_4 ( .A(puf_70_wire_0),  .B(puf_70_wire_6),  .S(sel), .Y(puf_70_wire_7));
   INVX1 puf_70_instance_5 ( .A(puf_70_wire_7), .Y(puf_70_wire_8));
   INVX1 puf_70_instance_6 ( .A(puf_70_wire_8), .Y(n85));
   BUFX2 puf_out_instance_70 ( .A(n85), .Y(pufout[70]));
   INVX1 puf_71_instance_0 ( .A(puf_71_wire_1), .Y(puf_71_wire_0));
   MUX2X1 puf_71_instance_1 ( .A(puf_71_wire_0),  .B(n86),  .S(sel), .Y(puf_71_wire_2));
   INVX1 puf_71_instance_2 ( .A(puf_71_wire_2), .Y(puf_71_wire_5));
   INVX1 puf_71_instance_3 ( .A(puf_71_wire_5), .Y(puf_71_wire_6));
   MUX2X1 puf_71_instance_4 ( .A(puf_71_wire_0),  .B(puf_71_wire_6),  .S(sel), .Y(puf_71_wire_7));
   INVX1 puf_71_instance_5 ( .A(puf_71_wire_7), .Y(puf_71_wire_8));
   INVX1 puf_71_instance_6 ( .A(puf_71_wire_8), .Y(n86));
   BUFX2 puf_out_instance_71 ( .A(n86), .Y(pufout[71]));
   INVX1 puf_72_instance_0 ( .A(puf_72_wire_1), .Y(puf_72_wire_0));
   MUX2X1 puf_72_instance_1 ( .A(puf_72_wire_0),  .B(n87),  .S(sel), .Y(puf_72_wire_2));
   INVX1 puf_72_instance_2 ( .A(puf_72_wire_2), .Y(puf_72_wire_5));
   INVX1 puf_72_instance_3 ( .A(puf_72_wire_5), .Y(puf_72_wire_6));
   MUX2X1 puf_72_instance_4 ( .A(puf_72_wire_0),  .B(puf_72_wire_6),  .S(sel), .Y(puf_72_wire_7));
   INVX1 puf_72_instance_5 ( .A(puf_72_wire_7), .Y(puf_72_wire_8));
   INVX1 puf_72_instance_6 ( .A(puf_72_wire_8), .Y(n87));
   BUFX2 puf_out_instance_72 ( .A(n87), .Y(pufout[72]));
   INVX1 puf_73_instance_0 ( .A(puf_73_wire_1), .Y(puf_73_wire_0));
   MUX2X1 puf_73_instance_1 ( .A(puf_73_wire_0),  .B(n88),  .S(sel), .Y(puf_73_wire_2));
   INVX1 puf_73_instance_2 ( .A(puf_73_wire_2), .Y(puf_73_wire_5));
   INVX1 puf_73_instance_3 ( .A(puf_73_wire_5), .Y(puf_73_wire_6));
   MUX2X1 puf_73_instance_4 ( .A(puf_73_wire_0),  .B(puf_73_wire_6),  .S(sel), .Y(puf_73_wire_7));
   INVX1 puf_73_instance_5 ( .A(puf_73_wire_7), .Y(puf_73_wire_8));
   INVX1 puf_73_instance_6 ( .A(puf_73_wire_8), .Y(n88));
   BUFX2 puf_out_instance_73 ( .A(n88), .Y(pufout[73]));
   INVX1 puf_74_instance_0 ( .A(puf_74_wire_1), .Y(puf_74_wire_0));
   MUX2X1 puf_74_instance_1 ( .A(puf_74_wire_0),  .B(n89),  .S(sel), .Y(puf_74_wire_2));
   INVX1 puf_74_instance_2 ( .A(puf_74_wire_2), .Y(puf_74_wire_5));
   INVX1 puf_74_instance_3 ( .A(puf_74_wire_5), .Y(puf_74_wire_6));
   MUX2X1 puf_74_instance_4 ( .A(puf_74_wire_0),  .B(puf_74_wire_6),  .S(sel), .Y(puf_74_wire_7));
   INVX1 puf_74_instance_5 ( .A(puf_74_wire_7), .Y(puf_74_wire_8));
   INVX1 puf_74_instance_6 ( .A(puf_74_wire_8), .Y(n89));
   BUFX2 puf_out_instance_74 ( .A(n89), .Y(pufout[74]));
   INVX1 puf_75_instance_0 ( .A(puf_75_wire_1), .Y(puf_75_wire_0));
   MUX2X1 puf_75_instance_1 ( .A(puf_75_wire_0),  .B(n90),  .S(sel), .Y(puf_75_wire_2));
   INVX1 puf_75_instance_2 ( .A(puf_75_wire_2), .Y(puf_75_wire_5));
   INVX1 puf_75_instance_3 ( .A(puf_75_wire_5), .Y(puf_75_wire_6));
   MUX2X1 puf_75_instance_4 ( .A(puf_75_wire_0),  .B(puf_75_wire_6),  .S(sel), .Y(puf_75_wire_7));
   INVX1 puf_75_instance_5 ( .A(puf_75_wire_7), .Y(puf_75_wire_8));
   INVX1 puf_75_instance_6 ( .A(puf_75_wire_8), .Y(n90));
   BUFX2 puf_out_instance_75 ( .A(n90), .Y(pufout[75]));
   INVX1 puf_76_instance_0 ( .A(puf_76_wire_1), .Y(puf_76_wire_0));
   MUX2X1 puf_76_instance_1 ( .A(puf_76_wire_0),  .B(n91),  .S(sel), .Y(puf_76_wire_2));
   INVX1 puf_76_instance_2 ( .A(puf_76_wire_2), .Y(puf_76_wire_5));
   INVX1 puf_76_instance_3 ( .A(puf_76_wire_5), .Y(puf_76_wire_6));
   MUX2X1 puf_76_instance_4 ( .A(puf_76_wire_0),  .B(puf_76_wire_6),  .S(sel), .Y(puf_76_wire_7));
   INVX1 puf_76_instance_5 ( .A(puf_76_wire_7), .Y(puf_76_wire_8));
   INVX1 puf_76_instance_6 ( .A(puf_76_wire_8), .Y(n91));
   BUFX2 puf_out_instance_76 ( .A(n91), .Y(pufout[76]));
   INVX1 puf_77_instance_0 ( .A(puf_77_wire_1), .Y(puf_77_wire_0));
   MUX2X1 puf_77_instance_1 ( .A(puf_77_wire_0),  .B(n92),  .S(sel), .Y(puf_77_wire_2));
   INVX1 puf_77_instance_2 ( .A(puf_77_wire_2), .Y(puf_77_wire_5));
   INVX1 puf_77_instance_3 ( .A(puf_77_wire_5), .Y(puf_77_wire_6));
   MUX2X1 puf_77_instance_4 ( .A(puf_77_wire_0),  .B(puf_77_wire_6),  .S(sel), .Y(puf_77_wire_7));
   INVX1 puf_77_instance_5 ( .A(puf_77_wire_7), .Y(puf_77_wire_8));
   INVX1 puf_77_instance_6 ( .A(puf_77_wire_8), .Y(n92));
   BUFX2 puf_out_instance_77 ( .A(n92), .Y(pufout[77]));
   INVX1 puf_78_instance_0 ( .A(puf_78_wire_1), .Y(puf_78_wire_0));
   MUX2X1 puf_78_instance_1 ( .A(puf_78_wire_0),  .B(n93),  .S(sel), .Y(puf_78_wire_2));
   INVX1 puf_78_instance_2 ( .A(puf_78_wire_2), .Y(puf_78_wire_5));
   INVX1 puf_78_instance_3 ( .A(puf_78_wire_5), .Y(puf_78_wire_6));
   MUX2X1 puf_78_instance_4 ( .A(puf_78_wire_0),  .B(puf_78_wire_6),  .S(sel), .Y(puf_78_wire_7));
   INVX1 puf_78_instance_5 ( .A(puf_78_wire_7), .Y(puf_78_wire_8));
   INVX1 puf_78_instance_6 ( .A(puf_78_wire_8), .Y(n93));
   BUFX2 puf_out_instance_78 ( .A(n93), .Y(pufout[78]));
   INVX1 puf_79_instance_0 ( .A(puf_79_wire_1), .Y(puf_79_wire_0));
   MUX2X1 puf_79_instance_1 ( .A(puf_79_wire_0),  .B(n94),  .S(sel), .Y(puf_79_wire_2));
   INVX1 puf_79_instance_2 ( .A(puf_79_wire_2), .Y(puf_79_wire_5));
   INVX1 puf_79_instance_3 ( .A(puf_79_wire_5), .Y(puf_79_wire_6));
   MUX2X1 puf_79_instance_4 ( .A(puf_79_wire_0),  .B(puf_79_wire_6),  .S(sel), .Y(puf_79_wire_7));
   INVX1 puf_79_instance_5 ( .A(puf_79_wire_7), .Y(puf_79_wire_8));
   INVX1 puf_79_instance_6 ( .A(puf_79_wire_8), .Y(n94));
   BUFX2 puf_out_instance_79 ( .A(n94), .Y(pufout[79]));
   INVX1 puf_80_instance_0 ( .A(puf_80_wire_1), .Y(puf_80_wire_0));
   MUX2X1 puf_80_instance_1 ( .A(puf_80_wire_0),  .B(n95),  .S(sel), .Y(puf_80_wire_2));
   INVX1 puf_80_instance_2 ( .A(puf_80_wire_2), .Y(puf_80_wire_5));
   INVX1 puf_80_instance_3 ( .A(puf_80_wire_5), .Y(puf_80_wire_6));
   MUX2X1 puf_80_instance_4 ( .A(puf_80_wire_0),  .B(puf_80_wire_6),  .S(sel), .Y(puf_80_wire_7));
   INVX1 puf_80_instance_5 ( .A(puf_80_wire_7), .Y(puf_80_wire_8));
   INVX1 puf_80_instance_6 ( .A(puf_80_wire_8), .Y(n95));
   BUFX2 puf_out_instance_80 ( .A(n95), .Y(pufout[80]));
   INVX1 puf_81_instance_0 ( .A(puf_81_wire_1), .Y(puf_81_wire_0));
   MUX2X1 puf_81_instance_1 ( .A(puf_81_wire_0),  .B(n96),  .S(sel), .Y(puf_81_wire_2));
   INVX1 puf_81_instance_2 ( .A(puf_81_wire_2), .Y(puf_81_wire_5));
   INVX1 puf_81_instance_3 ( .A(puf_81_wire_5), .Y(puf_81_wire_6));
   MUX2X1 puf_81_instance_4 ( .A(puf_81_wire_0),  .B(puf_81_wire_6),  .S(sel), .Y(puf_81_wire_7));
   INVX1 puf_81_instance_5 ( .A(puf_81_wire_7), .Y(puf_81_wire_8));
   INVX1 puf_81_instance_6 ( .A(puf_81_wire_8), .Y(n96));
   BUFX2 puf_out_instance_81 ( .A(n96), .Y(pufout[81]));
   INVX1 puf_82_instance_0 ( .A(puf_82_wire_1), .Y(puf_82_wire_0));
   MUX2X1 puf_82_instance_1 ( .A(puf_82_wire_0),  .B(n97),  .S(sel), .Y(puf_82_wire_2));
   INVX1 puf_82_instance_2 ( .A(puf_82_wire_2), .Y(puf_82_wire_5));
   INVX1 puf_82_instance_3 ( .A(puf_82_wire_5), .Y(puf_82_wire_6));
   MUX2X1 puf_82_instance_4 ( .A(puf_82_wire_0),  .B(puf_82_wire_6),  .S(sel), .Y(puf_82_wire_7));
   INVX1 puf_82_instance_5 ( .A(puf_82_wire_7), .Y(puf_82_wire_8));
   INVX1 puf_82_instance_6 ( .A(puf_82_wire_8), .Y(n97));
   BUFX2 puf_out_instance_82 ( .A(n97), .Y(pufout[82]));
   INVX1 puf_83_instance_0 ( .A(puf_83_wire_1), .Y(puf_83_wire_0));
   MUX2X1 puf_83_instance_1 ( .A(puf_83_wire_0),  .B(n98),  .S(sel), .Y(puf_83_wire_2));
   INVX1 puf_83_instance_2 ( .A(puf_83_wire_2), .Y(puf_83_wire_5));
   INVX1 puf_83_instance_3 ( .A(puf_83_wire_5), .Y(puf_83_wire_6));
   MUX2X1 puf_83_instance_4 ( .A(puf_83_wire_0),  .B(puf_83_wire_6),  .S(sel), .Y(puf_83_wire_7));
   INVX1 puf_83_instance_5 ( .A(puf_83_wire_7), .Y(puf_83_wire_8));
   INVX1 puf_83_instance_6 ( .A(puf_83_wire_8), .Y(n98));
   BUFX2 puf_out_instance_83 ( .A(n98), .Y(pufout[83]));
   INVX1 puf_84_instance_0 ( .A(puf_84_wire_1), .Y(puf_84_wire_0));
   MUX2X1 puf_84_instance_1 ( .A(puf_84_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[1]),  .S(sel), .Y(puf_84_wire_2));
   INVX1 puf_84_instance_2 ( .A(puf_84_wire_2), .Y(puf_84_wire_5));
   INVX1 puf_84_instance_3 ( .A(puf_84_wire_5), .Y(puf_84_wire_6));
   MUX2X1 puf_84_instance_4 ( .A(puf_84_wire_0),  .B(puf_84_wire_6),  .S(sel), .Y(puf_84_wire_7));
   INVX1 puf_84_instance_5 ( .A(puf_84_wire_7), .Y(puf_84_wire_8));
   INVX1 puf_84_instance_6 ( .A(puf_84_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[1]));
   BUFX2 puf_out_instance_84 ( .A(my_FIR_filter_firBlock_right_multProducts[1]), .Y(pufout[84]));
   INVX1 puf_85_instance_0 ( .A(puf_85_wire_1), .Y(puf_85_wire_0));
   MUX2X1 puf_85_instance_1 ( .A(puf_85_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[2]),  .S(sel), .Y(puf_85_wire_2));
   INVX1 puf_85_instance_2 ( .A(puf_85_wire_2), .Y(puf_85_wire_5));
   INVX1 puf_85_instance_3 ( .A(puf_85_wire_5), .Y(puf_85_wire_6));
   MUX2X1 puf_85_instance_4 ( .A(puf_85_wire_0),  .B(puf_85_wire_6),  .S(sel), .Y(puf_85_wire_7));
   INVX1 puf_85_instance_5 ( .A(puf_85_wire_7), .Y(puf_85_wire_8));
   INVX1 puf_85_instance_6 ( .A(puf_85_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[2]));
   BUFX2 puf_out_instance_85 ( .A(my_FIR_filter_firBlock_right_multProducts[2]), .Y(pufout[85]));
   INVX1 puf_86_instance_0 ( .A(puf_86_wire_1), .Y(puf_86_wire_0));
   MUX2X1 puf_86_instance_1 ( .A(puf_86_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[3]),  .S(sel), .Y(puf_86_wire_2));
   INVX1 puf_86_instance_2 ( .A(puf_86_wire_2), .Y(puf_86_wire_5));
   INVX1 puf_86_instance_3 ( .A(puf_86_wire_5), .Y(puf_86_wire_6));
   MUX2X1 puf_86_instance_4 ( .A(puf_86_wire_0),  .B(puf_86_wire_6),  .S(sel), .Y(puf_86_wire_7));
   INVX1 puf_86_instance_5 ( .A(puf_86_wire_7), .Y(puf_86_wire_8));
   INVX1 puf_86_instance_6 ( .A(puf_86_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[3]));
   BUFX2 puf_out_instance_86 ( .A(my_FIR_filter_firBlock_right_multProducts[3]), .Y(pufout[86]));
   INVX1 puf_87_instance_0 ( .A(puf_87_wire_1), .Y(puf_87_wire_0));
   MUX2X1 puf_87_instance_1 ( .A(puf_87_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[4]),  .S(sel), .Y(puf_87_wire_2));
   INVX1 puf_87_instance_2 ( .A(puf_87_wire_2), .Y(puf_87_wire_5));
   INVX1 puf_87_instance_3 ( .A(puf_87_wire_5), .Y(puf_87_wire_6));
   MUX2X1 puf_87_instance_4 ( .A(puf_87_wire_0),  .B(puf_87_wire_6),  .S(sel), .Y(puf_87_wire_7));
   INVX1 puf_87_instance_5 ( .A(puf_87_wire_7), .Y(puf_87_wire_8));
   INVX1 puf_87_instance_6 ( .A(puf_87_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[4]));
   BUFX2 puf_out_instance_87 ( .A(my_FIR_filter_firBlock_right_multProducts[4]), .Y(pufout[87]));
   INVX1 puf_88_instance_0 ( .A(puf_88_wire_1), .Y(puf_88_wire_0));
   MUX2X1 puf_88_instance_1 ( .A(puf_88_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[5]),  .S(sel), .Y(puf_88_wire_2));
   INVX1 puf_88_instance_2 ( .A(puf_88_wire_2), .Y(puf_88_wire_5));
   INVX1 puf_88_instance_3 ( .A(puf_88_wire_5), .Y(puf_88_wire_6));
   MUX2X1 puf_88_instance_4 ( .A(puf_88_wire_0),  .B(puf_88_wire_6),  .S(sel), .Y(puf_88_wire_7));
   INVX1 puf_88_instance_5 ( .A(puf_88_wire_7), .Y(puf_88_wire_8));
   INVX1 puf_88_instance_6 ( .A(puf_88_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[5]));
   BUFX2 puf_out_instance_88 ( .A(my_FIR_filter_firBlock_right_multProducts[5]), .Y(pufout[88]));
   INVX1 puf_89_instance_0 ( .A(puf_89_wire_1), .Y(puf_89_wire_0));
   MUX2X1 puf_89_instance_1 ( .A(puf_89_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[6]),  .S(sel), .Y(puf_89_wire_2));
   INVX1 puf_89_instance_2 ( .A(puf_89_wire_2), .Y(puf_89_wire_5));
   INVX1 puf_89_instance_3 ( .A(puf_89_wire_5), .Y(puf_89_wire_6));
   MUX2X1 puf_89_instance_4 ( .A(puf_89_wire_0),  .B(puf_89_wire_6),  .S(sel), .Y(puf_89_wire_7));
   INVX1 puf_89_instance_5 ( .A(puf_89_wire_7), .Y(puf_89_wire_8));
   INVX1 puf_89_instance_6 ( .A(puf_89_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[6]));
   BUFX2 puf_out_instance_89 ( .A(my_FIR_filter_firBlock_right_multProducts[6]), .Y(pufout[89]));
   INVX1 puf_90_instance_0 ( .A(puf_90_wire_1), .Y(puf_90_wire_0));
   MUX2X1 puf_90_instance_1 ( .A(puf_90_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[7]),  .S(sel), .Y(puf_90_wire_2));
   INVX1 puf_90_instance_2 ( .A(puf_90_wire_2), .Y(puf_90_wire_5));
   INVX1 puf_90_instance_3 ( .A(puf_90_wire_5), .Y(puf_90_wire_6));
   MUX2X1 puf_90_instance_4 ( .A(puf_90_wire_0),  .B(puf_90_wire_6),  .S(sel), .Y(puf_90_wire_7));
   INVX1 puf_90_instance_5 ( .A(puf_90_wire_7), .Y(puf_90_wire_8));
   INVX1 puf_90_instance_6 ( .A(puf_90_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[7]));
   BUFX2 puf_out_instance_90 ( .A(my_FIR_filter_firBlock_right_multProducts[7]), .Y(pufout[90]));
   INVX1 puf_91_instance_0 ( .A(puf_91_wire_1), .Y(puf_91_wire_0));
   MUX2X1 puf_91_instance_1 ( .A(puf_91_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[8]),  .S(sel), .Y(puf_91_wire_2));
   INVX1 puf_91_instance_2 ( .A(puf_91_wire_2), .Y(puf_91_wire_5));
   INVX1 puf_91_instance_3 ( .A(puf_91_wire_5), .Y(puf_91_wire_6));
   MUX2X1 puf_91_instance_4 ( .A(puf_91_wire_0),  .B(puf_91_wire_6),  .S(sel), .Y(puf_91_wire_7));
   INVX1 puf_91_instance_5 ( .A(puf_91_wire_7), .Y(puf_91_wire_8));
   INVX1 puf_91_instance_6 ( .A(puf_91_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[8]));
   BUFX2 puf_out_instance_91 ( .A(my_FIR_filter_firBlock_right_multProducts[8]), .Y(pufout[91]));
   INVX1 puf_92_instance_0 ( .A(puf_92_wire_1), .Y(puf_92_wire_0));
   MUX2X1 puf_92_instance_1 ( .A(puf_92_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[9]),  .S(sel), .Y(puf_92_wire_2));
   INVX1 puf_92_instance_2 ( .A(puf_92_wire_2), .Y(puf_92_wire_5));
   INVX1 puf_92_instance_3 ( .A(puf_92_wire_5), .Y(puf_92_wire_6));
   MUX2X1 puf_92_instance_4 ( .A(puf_92_wire_0),  .B(puf_92_wire_6),  .S(sel), .Y(puf_92_wire_7));
   INVX1 puf_92_instance_5 ( .A(puf_92_wire_7), .Y(puf_92_wire_8));
   INVX1 puf_92_instance_6 ( .A(puf_92_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[9]));
   BUFX2 puf_out_instance_92 ( .A(my_FIR_filter_firBlock_right_multProducts[9]), .Y(pufout[92]));
   INVX1 puf_93_instance_0 ( .A(puf_93_wire_1), .Y(puf_93_wire_0));
   MUX2X1 puf_93_instance_1 ( .A(puf_93_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[10]),  .S(sel), .Y(puf_93_wire_2));
   INVX1 puf_93_instance_2 ( .A(puf_93_wire_2), .Y(puf_93_wire_5));
   INVX1 puf_93_instance_3 ( .A(puf_93_wire_5), .Y(puf_93_wire_6));
   MUX2X1 puf_93_instance_4 ( .A(puf_93_wire_0),  .B(puf_93_wire_6),  .S(sel), .Y(puf_93_wire_7));
   INVX1 puf_93_instance_5 ( .A(puf_93_wire_7), .Y(puf_93_wire_8));
   INVX1 puf_93_instance_6 ( .A(puf_93_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[10]));
   BUFX2 puf_out_instance_93 ( .A(my_FIR_filter_firBlock_right_multProducts[10]), .Y(pufout[93]));
   INVX1 puf_94_instance_0 ( .A(puf_94_wire_1), .Y(puf_94_wire_0));
   MUX2X1 puf_94_instance_1 ( .A(puf_94_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[11]),  .S(sel), .Y(puf_94_wire_2));
   INVX1 puf_94_instance_2 ( .A(puf_94_wire_2), .Y(puf_94_wire_5));
   INVX1 puf_94_instance_3 ( .A(puf_94_wire_5), .Y(puf_94_wire_6));
   MUX2X1 puf_94_instance_4 ( .A(puf_94_wire_0),  .B(puf_94_wire_6),  .S(sel), .Y(puf_94_wire_7));
   INVX1 puf_94_instance_5 ( .A(puf_94_wire_7), .Y(puf_94_wire_8));
   INVX1 puf_94_instance_6 ( .A(puf_94_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[11]));
   BUFX2 puf_out_instance_94 ( .A(my_FIR_filter_firBlock_right_multProducts[11]), .Y(pufout[94]));
   INVX1 puf_95_instance_0 ( .A(puf_95_wire_1), .Y(puf_95_wire_0));
   MUX2X1 puf_95_instance_1 ( .A(puf_95_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[12]),  .S(sel), .Y(puf_95_wire_2));
   INVX1 puf_95_instance_2 ( .A(puf_95_wire_2), .Y(puf_95_wire_5));
   INVX1 puf_95_instance_3 ( .A(puf_95_wire_5), .Y(puf_95_wire_6));
   MUX2X1 puf_95_instance_4 ( .A(puf_95_wire_0),  .B(puf_95_wire_6),  .S(sel), .Y(puf_95_wire_7));
   INVX1 puf_95_instance_5 ( .A(puf_95_wire_7), .Y(puf_95_wire_8));
   INVX1 puf_95_instance_6 ( .A(puf_95_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[12]));
   BUFX2 puf_out_instance_95 ( .A(my_FIR_filter_firBlock_right_multProducts[12]), .Y(pufout[95]));
   INVX1 puf_96_instance_0 ( .A(puf_96_wire_1), .Y(puf_96_wire_0));
   MUX2X1 puf_96_instance_1 ( .A(puf_96_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[13]),  .S(sel), .Y(puf_96_wire_2));
   INVX1 puf_96_instance_2 ( .A(puf_96_wire_2), .Y(puf_96_wire_5));
   INVX1 puf_96_instance_3 ( .A(puf_96_wire_5), .Y(puf_96_wire_6));
   MUX2X1 puf_96_instance_4 ( .A(puf_96_wire_0),  .B(puf_96_wire_6),  .S(sel), .Y(puf_96_wire_7));
   INVX1 puf_96_instance_5 ( .A(puf_96_wire_7), .Y(puf_96_wire_8));
   INVX1 puf_96_instance_6 ( .A(puf_96_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[13]));
   BUFX2 puf_out_instance_96 ( .A(my_FIR_filter_firBlock_right_multProducts[13]), .Y(pufout[96]));
   INVX1 puf_97_instance_0 ( .A(puf_97_wire_1), .Y(puf_97_wire_0));
   MUX2X1 puf_97_instance_1 ( .A(puf_97_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[14]),  .S(sel), .Y(puf_97_wire_2));
   INVX1 puf_97_instance_2 ( .A(puf_97_wire_2), .Y(puf_97_wire_5));
   INVX1 puf_97_instance_3 ( .A(puf_97_wire_5), .Y(puf_97_wire_6));
   MUX2X1 puf_97_instance_4 ( .A(puf_97_wire_0),  .B(puf_97_wire_6),  .S(sel), .Y(puf_97_wire_7));
   INVX1 puf_97_instance_5 ( .A(puf_97_wire_7), .Y(puf_97_wire_8));
   INVX1 puf_97_instance_6 ( .A(puf_97_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[14]));
   BUFX2 puf_out_instance_97 ( .A(my_FIR_filter_firBlock_right_multProducts[14]), .Y(pufout[97]));
   INVX1 puf_98_instance_0 ( .A(puf_98_wire_1), .Y(puf_98_wire_0));
   MUX2X1 puf_98_instance_1 ( .A(puf_98_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[15]),  .S(sel), .Y(puf_98_wire_2));
   INVX1 puf_98_instance_2 ( .A(puf_98_wire_2), .Y(puf_98_wire_5));
   INVX1 puf_98_instance_3 ( .A(puf_98_wire_5), .Y(puf_98_wire_6));
   MUX2X1 puf_98_instance_4 ( .A(puf_98_wire_0),  .B(puf_98_wire_6),  .S(sel), .Y(puf_98_wire_7));
   INVX1 puf_98_instance_5 ( .A(puf_98_wire_7), .Y(puf_98_wire_8));
   INVX1 puf_98_instance_6 ( .A(puf_98_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[15]));
   BUFX2 puf_out_instance_98 ( .A(my_FIR_filter_firBlock_right_multProducts[15]), .Y(pufout[98]));
   INVX1 puf_99_instance_0 ( .A(puf_99_wire_1), .Y(puf_99_wire_0));
   MUX2X1 puf_99_instance_1 ( .A(puf_99_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[16]),  .S(sel), .Y(puf_99_wire_2));
   INVX1 puf_99_instance_2 ( .A(puf_99_wire_2), .Y(puf_99_wire_5));
   INVX1 puf_99_instance_3 ( .A(puf_99_wire_5), .Y(puf_99_wire_6));
   MUX2X1 puf_99_instance_4 ( .A(puf_99_wire_0),  .B(puf_99_wire_6),  .S(sel), .Y(puf_99_wire_7));
   INVX1 puf_99_instance_5 ( .A(puf_99_wire_7), .Y(puf_99_wire_8));
   INVX1 puf_99_instance_6 ( .A(puf_99_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[16]));
   BUFX2 puf_out_instance_99 ( .A(my_FIR_filter_firBlock_right_multProducts[16]), .Y(pufout[99]));
   INVX1 puf_100_instance_0 ( .A(puf_100_wire_1), .Y(puf_100_wire_0));
   MUX2X1 puf_100_instance_1 ( .A(puf_100_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[17]),  .S(sel), .Y(puf_100_wire_2));
   INVX1 puf_100_instance_2 ( .A(puf_100_wire_2), .Y(puf_100_wire_5));
   INVX1 puf_100_instance_3 ( .A(puf_100_wire_5), .Y(puf_100_wire_6));
   MUX2X1 puf_100_instance_4 ( .A(puf_100_wire_0),  .B(puf_100_wire_6),  .S(sel), .Y(puf_100_wire_7));
   INVX1 puf_100_instance_5 ( .A(puf_100_wire_7), .Y(puf_100_wire_8));
   INVX1 puf_100_instance_6 ( .A(puf_100_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[17]));
   BUFX2 puf_out_instance_100 ( .A(my_FIR_filter_firBlock_right_multProducts[17]), .Y(pufout[100]));
   INVX1 puf_101_instance_0 ( .A(puf_101_wire_1), .Y(puf_101_wire_0));
   MUX2X1 puf_101_instance_1 ( .A(puf_101_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[18]),  .S(sel), .Y(puf_101_wire_2));
   INVX1 puf_101_instance_2 ( .A(puf_101_wire_2), .Y(puf_101_wire_5));
   INVX1 puf_101_instance_3 ( .A(puf_101_wire_5), .Y(puf_101_wire_6));
   MUX2X1 puf_101_instance_4 ( .A(puf_101_wire_0),  .B(puf_101_wire_6),  .S(sel), .Y(puf_101_wire_7));
   INVX1 puf_101_instance_5 ( .A(puf_101_wire_7), .Y(puf_101_wire_8));
   INVX1 puf_101_instance_6 ( .A(puf_101_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[18]));
   BUFX2 puf_out_instance_101 ( .A(my_FIR_filter_firBlock_right_multProducts[18]), .Y(pufout[101]));
   INVX1 puf_102_instance_0 ( .A(puf_102_wire_1), .Y(puf_102_wire_0));
   MUX2X1 puf_102_instance_1 ( .A(puf_102_wire_0),  .B(my_FIR_filter_firBlock_right_multProducts[19]),  .S(sel), .Y(puf_102_wire_2));
   INVX1 puf_102_instance_2 ( .A(puf_102_wire_2), .Y(puf_102_wire_5));
   INVX1 puf_102_instance_3 ( .A(puf_102_wire_5), .Y(puf_102_wire_6));
   MUX2X1 puf_102_instance_4 ( .A(puf_102_wire_0),  .B(puf_102_wire_6),  .S(sel), .Y(puf_102_wire_7));
   INVX1 puf_102_instance_5 ( .A(puf_102_wire_7), .Y(puf_102_wire_8));
   INVX1 puf_102_instance_6 ( .A(puf_102_wire_8), .Y(my_FIR_filter_firBlock_right_multProducts[19]));
   BUFX2 puf_out_instance_102 ( .A(my_FIR_filter_firBlock_right_multProducts[19]), .Y(pufout[102]));
   INVX1 puf_103_instance_0 ( .A(puf_103_wire_1), .Y(puf_103_wire_0));
   MUX2X1 puf_103_instance_1 ( .A(puf_103_wire_0),  .B(my_FIR_filter_firBlock_left_N1),  .S(sel), .Y(puf_103_wire_2));
   INVX1 puf_103_instance_2 ( .A(puf_103_wire_2), .Y(puf_103_wire_5));
   INVX1 puf_103_instance_3 ( .A(puf_103_wire_5), .Y(puf_103_wire_6));
   MUX2X1 puf_103_instance_4 ( .A(puf_103_wire_0),  .B(puf_103_wire_6),  .S(sel), .Y(puf_103_wire_7));
   INVX1 puf_103_instance_5 ( .A(puf_103_wire_7), .Y(puf_103_wire_8));
   INVX1 puf_103_instance_6 ( .A(puf_103_wire_8), .Y(my_FIR_filter_firBlock_left_N1));
   BUFX2 puf_out_instance_103 ( .A(my_FIR_filter_firBlock_left_N1), .Y(pufout[103]));
   INVX1 puf_104_instance_0 ( .A(puf_104_wire_1), .Y(puf_104_wire_0));
   MUX2X1 puf_104_instance_1 ( .A(puf_104_wire_0),  .B(my_FIR_filter_firBlock_left_N33),  .S(sel), .Y(puf_104_wire_2));
   INVX1 puf_104_instance_2 ( .A(puf_104_wire_2), .Y(puf_104_wire_5));
   INVX1 puf_104_instance_3 ( .A(puf_104_wire_5), .Y(puf_104_wire_6));
   MUX2X1 puf_104_instance_4 ( .A(puf_104_wire_0),  .B(puf_104_wire_6),  .S(sel), .Y(puf_104_wire_7));
   INVX1 puf_104_instance_5 ( .A(puf_104_wire_7), .Y(puf_104_wire_8));
   INVX1 puf_104_instance_6 ( .A(puf_104_wire_8), .Y(my_FIR_filter_firBlock_left_N33));
   BUFX2 puf_out_instance_104 ( .A(my_FIR_filter_firBlock_left_N33), .Y(pufout[104]));
   INVX1 puf_105_instance_0 ( .A(puf_105_wire_1), .Y(puf_105_wire_0));
   MUX2X1 puf_105_instance_1 ( .A(puf_105_wire_0),  .B(my_FIR_filter_firBlock_left_N65),  .S(sel), .Y(puf_105_wire_2));
   INVX1 puf_105_instance_2 ( .A(puf_105_wire_2), .Y(puf_105_wire_5));
   INVX1 puf_105_instance_3 ( .A(puf_105_wire_5), .Y(puf_105_wire_6));
   MUX2X1 puf_105_instance_4 ( .A(puf_105_wire_0),  .B(puf_105_wire_6),  .S(sel), .Y(puf_105_wire_7));
   INVX1 puf_105_instance_5 ( .A(puf_105_wire_7), .Y(puf_105_wire_8));
   INVX1 puf_105_instance_6 ( .A(puf_105_wire_8), .Y(my_FIR_filter_firBlock_left_N65));
   BUFX2 puf_out_instance_105 ( .A(my_FIR_filter_firBlock_left_N65), .Y(pufout[105]));
   INVX1 puf_106_instance_0 ( .A(puf_106_wire_1), .Y(puf_106_wire_0));
   MUX2X1 puf_106_instance_1 ( .A(puf_106_wire_0),  .B(my_FIR_filter_firBlock_left_N97),  .S(sel), .Y(puf_106_wire_2));
   INVX1 puf_106_instance_2 ( .A(puf_106_wire_2), .Y(puf_106_wire_5));
   INVX1 puf_106_instance_3 ( .A(puf_106_wire_5), .Y(puf_106_wire_6));
   MUX2X1 puf_106_instance_4 ( .A(puf_106_wire_0),  .B(puf_106_wire_6),  .S(sel), .Y(puf_106_wire_7));
   INVX1 puf_106_instance_5 ( .A(puf_106_wire_7), .Y(puf_106_wire_8));
   INVX1 puf_106_instance_6 ( .A(puf_106_wire_8), .Y(my_FIR_filter_firBlock_left_N97));
   BUFX2 puf_out_instance_106 ( .A(my_FIR_filter_firBlock_left_N97), .Y(pufout[106]));
   INVX1 puf_107_instance_0 ( .A(puf_107_wire_1), .Y(puf_107_wire_0));
   MUX2X1 puf_107_instance_1 ( .A(puf_107_wire_0),  .B(my_FIR_filter_firBlock_left_N129),  .S(sel), .Y(puf_107_wire_2));
   INVX1 puf_107_instance_2 ( .A(puf_107_wire_2), .Y(puf_107_wire_5));
   INVX1 puf_107_instance_3 ( .A(puf_107_wire_5), .Y(puf_107_wire_6));
   MUX2X1 puf_107_instance_4 ( .A(puf_107_wire_0),  .B(puf_107_wire_6),  .S(sel), .Y(puf_107_wire_7));
   INVX1 puf_107_instance_5 ( .A(puf_107_wire_7), .Y(puf_107_wire_8));
   INVX1 puf_107_instance_6 ( .A(puf_107_wire_8), .Y(my_FIR_filter_firBlock_left_N129));
   BUFX2 puf_out_instance_107 ( .A(my_FIR_filter_firBlock_left_N129), .Y(pufout[107]));
   INVX1 puf_108_instance_0 ( .A(puf_108_wire_1), .Y(puf_108_wire_0));
   MUX2X1 puf_108_instance_1 ( .A(puf_108_wire_0),  .B(my_FIR_filter_firBlock_left_N161),  .S(sel), .Y(puf_108_wire_2));
   INVX1 puf_108_instance_2 ( .A(puf_108_wire_2), .Y(puf_108_wire_5));
   INVX1 puf_108_instance_3 ( .A(puf_108_wire_5), .Y(puf_108_wire_6));
   MUX2X1 puf_108_instance_4 ( .A(puf_108_wire_0),  .B(puf_108_wire_6),  .S(sel), .Y(puf_108_wire_7));
   INVX1 puf_108_instance_5 ( .A(puf_108_wire_7), .Y(puf_108_wire_8));
   INVX1 puf_108_instance_6 ( .A(puf_108_wire_8), .Y(my_FIR_filter_firBlock_left_N161));
   BUFX2 puf_out_instance_108 ( .A(my_FIR_filter_firBlock_left_N161), .Y(pufout[108]));
   INVX1 puf_109_instance_0 ( .A(puf_109_wire_1), .Y(puf_109_wire_0));
   MUX2X1 puf_109_instance_1 ( .A(puf_109_wire_0),  .B(my_FIR_filter_firBlock_left_N193),  .S(sel), .Y(puf_109_wire_2));
   INVX1 puf_109_instance_2 ( .A(puf_109_wire_2), .Y(puf_109_wire_5));
   INVX1 puf_109_instance_3 ( .A(puf_109_wire_5), .Y(puf_109_wire_6));
   MUX2X1 puf_109_instance_4 ( .A(puf_109_wire_0),  .B(puf_109_wire_6),  .S(sel), .Y(puf_109_wire_7));
   INVX1 puf_109_instance_5 ( .A(puf_109_wire_7), .Y(puf_109_wire_8));
   INVX1 puf_109_instance_6 ( .A(puf_109_wire_8), .Y(my_FIR_filter_firBlock_left_N193));
   BUFX2 puf_out_instance_109 ( .A(my_FIR_filter_firBlock_left_N193), .Y(pufout[109]));
   INVX1 puf_110_instance_0 ( .A(puf_110_wire_1), .Y(puf_110_wire_0));
   MUX2X1 puf_110_instance_1 ( .A(puf_110_wire_0),  .B(my_FIR_filter_firBlock_left_N225),  .S(sel), .Y(puf_110_wire_2));
   INVX1 puf_110_instance_2 ( .A(puf_110_wire_2), .Y(puf_110_wire_5));
   INVX1 puf_110_instance_3 ( .A(puf_110_wire_5), .Y(puf_110_wire_6));
   MUX2X1 puf_110_instance_4 ( .A(puf_110_wire_0),  .B(puf_110_wire_6),  .S(sel), .Y(puf_110_wire_7));
   INVX1 puf_110_instance_5 ( .A(puf_110_wire_7), .Y(puf_110_wire_8));
   INVX1 puf_110_instance_6 ( .A(puf_110_wire_8), .Y(my_FIR_filter_firBlock_left_N225));
   BUFX2 puf_out_instance_110 ( .A(my_FIR_filter_firBlock_left_N225), .Y(pufout[110]));
   INVX1 puf_111_instance_0 ( .A(puf_111_wire_1), .Y(puf_111_wire_0));
   MUX2X1 puf_111_instance_1 ( .A(puf_111_wire_0),  .B(my_FIR_filter_firBlock_left_N257),  .S(sel), .Y(puf_111_wire_2));
   INVX1 puf_111_instance_2 ( .A(puf_111_wire_2), .Y(puf_111_wire_5));
   INVX1 puf_111_instance_3 ( .A(puf_111_wire_5), .Y(puf_111_wire_6));
   MUX2X1 puf_111_instance_4 ( .A(puf_111_wire_0),  .B(puf_111_wire_6),  .S(sel), .Y(puf_111_wire_7));
   INVX1 puf_111_instance_5 ( .A(puf_111_wire_7), .Y(puf_111_wire_8));
   INVX1 puf_111_instance_6 ( .A(puf_111_wire_8), .Y(my_FIR_filter_firBlock_left_N257));
   BUFX2 puf_out_instance_111 ( .A(my_FIR_filter_firBlock_left_N257), .Y(pufout[111]));
endmodule


