.SUBCKT ad INOUT
M1 AIO VSS VSS VSS nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and2s1 Q DIN1 DIN2
M1 N1N251 DIN1 VDD VDD pch W=0.7U L=0.24U
M2 N1N251 DIN2 VDD VDD pch W=0.7U L=0.24U
M3 N1N251 DIN1 N1N257 VSS nch W=0.7U L=0.24U
M4 N1N257 DIN2 VSS VSS nch W=0.7U L=0.24U
M5 Q N1N251 VDD VDD pch W=1.76U L=0.24U
M6 Q N1N251 VSS VSS nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and2s2 Q DIN1 DIN2
M3 N1N257 DIN1 N1N259 VSS nch W=2.14U L=0.24U
M1 N1N257 DIN1 VDD VDD pch W=2.4U L=0.24U
M2 N1N257 DIN2 VDD VDD pch W=2.4U L=0.24U
M5 Q N1N257 VDD VDD pch W=5.3U L=0.24U
M4 N1N259 DIN2 VSS VSS nch W=2.14U L=0.24U
M6 Q N1N257 VSS VSS nch W=3.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and2s3 Q DIN1 DIN2
M3 N1N257 DIN1 N1N259 VSS nch W=4.4U L=0.24U
M1 N1N257 DIN1 VDD VDD pch W=4.5U L=0.24U
M2 N1N257 DIN2 VDD VDD pch W=4.5U L=0.24U
M4 N1N259 DIN2 VSS VSS nch W=4.4U L=0.24U
M5 Q N1N257 VDD VDD pch W=9.5U L=0.24U
M6 Q N1N257 VSS VSS nch W=6.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and3s1 Q DIN1 DIN2 DIN3
M4 N1N258 DIN1 N1N262 VSS nch W=1.08U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=0.82U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=0.82U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=0.82U L=0.24U
M5 N1N262 DIN2 N1N264 VSS nch W=1.08U L=0.24U
M6 N1N264 DIN3 VSS VSS nch W=1.08U L=0.24U
M8 Q N1N258 VSS VSS nch W=1.34U L=0.24U
M7 Q N1N258 VDD VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and3s2 Q DIN1 DIN2 DIN3
M4 N1N258 DIN1 N1N262 VSS nch W=3.14U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=2.54U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=2.54U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=2.54U L=0.24U
M5 N1N262 DIN2 N1N264 VSS nch W=3.14U L=0.24U
M6 N1N264 DIN3 VSS VSS nch W=3.14U L=0.24U
M8 Q N1N258 VSS VSS nch W=4.1U L=0.24U
M7 Q N1N258 VDD VDD pch W=4.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and3s3 Q DIN1 DIN2 DIN3
M4 N1N258 DIN1 N1N262 VSS nch W=3.8U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=4.7U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=4.7U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=4.7U L=0.24U
M5 N1N262 DIN2 N1N264 VSS nch W=4.76U L=0.24U
M6 N1N264 DIN3 VSS VSS nch W=7.4U L=0.24U
M8 Q N1N258 VSS VSS nch W=7.4U L=0.24U
M7 Q N1N258 VDD VDD pch W=9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and4s1 Q DIN1 DIN2 DIN3 DIN4
M5 N1N258 DIN1 N1N265 VSS nch W=1U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=1U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=1U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=1U L=0.24U
M4 N1N258 DIN4 VDD VDD pch W=1U L=0.24U
M6 N1N265 DIN2 N1N267 VSS nch W=1.24U L=0.24U
M7 N1N267 DIN3 N1N269 VSS nch W=1.44U L=0.24U
M8 N1N269 DIN4 VSS VSS nch W=1.64U L=0.24U
M9 Q N1N258 VDD VDD pch W=1.96U L=0.24U
M10 Q N1N258 VSS VSS nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and4s2 Q DIN1 DIN2 DIN3 DIN4
M5 N1N258 DIN1 N1N265 VSS nch W=2.32U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=3U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=3U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=3U L=0.24U
M4 N1N258 DIN4 VDD VDD pch W=3U L=0.24U
M6 N1N265 DIN2 N1N267 VSS nch W=2.54U L=0.24U
M7 N1N267 DIN3 N1N269 VSS nch W=3.96U L=0.24U
M8 N1N269 DIN4 VSS VSS nch W=4.16U L=0.24U
M9 Q N1N258 VDD VDD pch W=5.7U L=0.24U
M10 Q N1N258 VSS VSS nch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and4s3 DIN1 DIN2 DIN3 DIN4 Q
M3 N1N259 DIN1 N1N262 VSS nch W=3.16U L=0.24U
M1 N1N259 DIN1 VDD VDD pch W=3.5U L=0.24U
M2 VDD DIN2 N1N259 VDD pch W=3.5U L=0.24U
M4 N1N262 DIN2 VSS VSS nch W=4.1U L=0.24U
M9 N1N279 N1N259 VDD VDD pch W=7.2U L=0.24U
M10 N1N279 N1N270 Q VDD pch W=7U L=0.24U
M5 N1N270 DIN3 VDD VDD pch W=3.5U L=0.24U
M6 VDD DIN4 N1N270 VDD pch W=3.5U L=0.24U
M7 N1N270 DIN3 N1N273 VSS nch W=3.16U L=0.24U
M8 N1N273 DIN4 VSS VSS nch W=4.1U L=0.24U
M11 Q N1N259 VSS VSS nch W=2.5U L=0.24U
M12 VSS N1N270 Q VSS nch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoai1112s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N286 DIN1 Q VSS nch W=0.8U L=0.24U
M1 N1N282 DIN4 VDD VDD pch W=1.5U L=0.24U
M2 N1N282 DIN5 VDD VDD pch W=1.5U L=0.24U
M3 Q DIN3 N1N282 VDD pch W=1.4U L=0.24U
M4 VDD DIN2 Q VDD pch W=0.7U L=0.24U
M5 VDD DIN1 Q VDD pch W=0.7U L=0.24U
M7 N1N299 DIN2 N1N286 VSS nch W=0.8U L=0.24U
M8 N1N299 DIN3 VSS VSS nch W=0.8U L=0.24U
M9 N1N299 DIN4 N1N302 VSS nch W=1.6U L=0.24U
M10 N1N302 DIN5 VSS VSS nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoai1112s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N286 DIN1 Q VSS nch W=1.1U L=0.24U
M1 N1N282 DIN4 VDD VDD pch W=2U L=0.24U
M2 N1N282 DIN5 VDD VDD pch W=2U L=0.24U
M3 Q DIN3 N1N282 VDD pch W=1.9U L=0.24U
M4 VDD DIN2 Q VDD pch W=1U L=0.24U
M5 VDD DIN1 Q VDD pch W=1U L=0.24U
M7 N1N299 DIN2 N1N286 VSS nch W=1.1U L=0.24U
M8 N1N299 DIN3 VSS VSS nch W=1.1U L=0.24U
M9 N1N299 DIN4 N1N302 VSS nch W=2.2U L=0.24U
M10 N1N302 DIN5 VSS VSS nch W=2.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoai1112s3 DIN1 DIN2 DIN3 DIN4 DIN5 Q
M6 N1N286 DIN1 Q VSS nch W=1.6U L=0.24U
M1 N1N282 DIN4 VDD VDD pch W=3.3U L=0.24U
M2 N1N282 DIN5 VDD VDD pch W=3.4U L=0.24U
M3 Q DIN3 N1N282 VDD pch W=3.3U L=0.24U
M4 VDD DIN2 Q VDD pch W=1.7U L=0.24U
M5 VDD DIN1 Q VDD pch W=1.7U L=0.24U
M7 N1N299 DIN2 N1N286 VSS nch W=1.7U L=0.24U
M8 N1N299 DIN3 VSS VSS nch W=1.7U L=0.24U
M9 N1N299 DIN4 N1N302 VSS nch W=3.4U L=0.24U
M10 N1N302 DIN5 VSS VSS nch W=3.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoai122s1 DIN1 DIN2 DIN3 DIN4 DIN5 Q
M6 Q DIN1 N1N298 VSS nch W=0.9U L=0.24U
M2 N1N290 DIN2 VDD VDD pch W=1.5U L=0.24U
M3 Q DIN4 N1N290 VDD pch W=1.5U L=0.24U
M4 VDD DIN3 N1N290 VDD pch W=1.5U L=0.24U
M5 N1N290 DIN5 Q VDD pch W=1.5U L=0.24U
M7 N1N298 DIN2 N1N300 VSS nch W=0.9U L=0.24U
M10 VSS DIN5 N1N302 VSS nch W=0.9U L=0.24U
M9 N1N302 DIN4 N1N298 VSS nch W=0.9U L=0.24U
M8 VSS DIN3 N1N300 VSS nch W=0.9U L=0.24U
M1 Q DIN1 VDD VDD pch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoai122s2 DIN1 DIN2 DIN3 DIN4 DIN5 Q
M6 Q DIN1 N1N298 VSS nch W=1.1U L=0.24U
M2 N1N290 DIN2 VDD VDD pch W=1.8U L=0.24U
M3 Q DIN4 N1N290 VDD pch W=1.8U L=0.24U
M4 VDD DIN3 N1N290 VDD pch W=1.8U L=0.24U
M5 N1N290 DIN5 Q VDD pch W=1.8U L=0.24U
M7 N1N298 DIN2 N1N300 VSS nch W=1.1U L=0.24U
M10 VSS DIN5 N1N302 VSS nch W=1.1U L=0.24U
M9 N1N302 DIN4 N1N298 VSS nch W=1.1U L=0.24U
M8 VSS DIN3 N1N300 VSS nch W=1.1U L=0.24U
M1 Q DIN1 VDD VDD pch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoai122s3 DIN1 DIN2 DIN3 DIN4 DIN5 Q
M6 N1N292 DIN1 N1N298 VSS nch W=0.9U L=0.24U
M2 N1N290 DIN2 VDD VDD pch W=1.5U L=0.24U
M3 N1N292 DIN4 N1N290 VDD pch W=1.5U L=0.24U
M4 VDD DIN3 N1N290 VDD pch W=1.5U L=0.24U
M5 N1N290 DIN5 N1N292 VDD pch W=1.5U L=0.24U
M7 N1N298 DIN2 N1N300 VSS nch W=1U L=0.24U
M10 VSS DIN5 N1N302 VSS nch W=1U L=0.24U
M9 N1N302 DIN4 N1N298 VSS nch W=1U L=0.24U
M8 VSS DIN3 N1N300 VSS nch W=1U L=0.24U
M1 N1N292 DIN1 VDD VDD pch W=0.7U L=0.24U
M12 N1N339 N1N292 VSS VSS nch W=1.4U L=0.24U
M11 N1N339 N1N292 VDD VDD pch W=2.7U L=0.24U
M13 Q N1N339 VDD VDD pch W=4.5U L=0.24U
M14 Q N1N339 VSS VSS nch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi123s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N461 DIN3 N1N445 VDD pch W=4.1U L=0.24U
M1 N1N445 DIN5 VDD VDD pch W=4.1U L=0.24U
M2 VDD DIN4 N1N445 VDD pch W=4.1U L=0.24U
M3 VDD DIN6 N1N445 VDD pch W=4.1U L=0.24U
M5 N1N445 DIN2 N1N461 VDD pch W=4.1U L=0.24U
M6 Q DIN1 N1N461 VDD pch W=4.1U L=0.24U
M7 N1N469 DIN2 Q VSS nch W=1.2U L=0.24U
M10 N1N469 DIN3 VSS VSS nch W=1.2U L=0.24U
M8 N1N473 DIN4 Q VSS nch W=1.8U L=0.24U
M12 VSS DIN6 N1N475 VSS nch W=1.8U L=0.24U
M11 N1N475 DIN5 N1N473 VSS nch W=1.8U L=0.24U
M9 Q DIN1 VSS VSS nch W=0.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi123s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N461 DIN3 N1N445 VDD pch W=5.8U L=0.24U
M1 N1N445 DIN5 VDD VDD pch W=5.8U L=0.24U
M2 VDD DIN4 N1N445 VDD pch W=5.8U L=0.24U
M3 VDD DIN6 N1N445 VDD pch W=5.8U L=0.24U
M5 N1N445 DIN2 N1N461 VDD pch W=5.8U L=0.24U
M6 Q DIN1 N1N461 VDD pch W=5.8U L=0.24U
M7 N1N469 DIN2 Q VSS nch W=1.7U L=0.24U
M10 N1N469 DIN3 VSS VSS nch W=1.7U L=0.24U
M8 N1N473 DIN4 Q VSS nch W=2.5U L=0.24U
M12 VSS DIN6 N1N475 VSS nch W=2.5U L=0.24U
M11 N1N475 DIN5 N1N473 VSS nch W=2.5U L=0.24U
M9 Q DIN1 VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi123s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N461 DIN3 N1N445 VDD pch W=7.8U L=0.24U
M1 N1N445 DIN5 VDD VDD pch W=7.8U L=0.24U
M2 VDD DIN4 N1N445 VDD pch W=7.8U L=0.24U
M3 VDD DIN6 N1N445 VDD pch W=7.8U L=0.24U
M5 N1N445 DIN2 N1N461 VDD pch W=7.8U L=0.24U
M6 Q DIN1 N1N461 VDD pch W=7.8U L=0.24U
M7 N1N469 DIN2 Q VSS nch W=2.2U L=0.24U
M10 N1N469 DIN3 VSS VSS nch W=2.2U L=0.24U
M8 N1N473 DIN4 Q VSS nch W=3.3U L=0.24U
M12 VSS DIN6 N1N475 VSS nch W=3.3U L=0.24U
M11 N1N475 DIN5 N1N473 VSS nch W=3.3U L=0.24U
M9 Q DIN1 VSS VSS nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi13s1 Q DIN1 DIN2 DIN3 DIN4
M6 N1N452 DIN2 Q VSS nch W=1.24U L=0.24U
M2 VDD DIN3 N1N490 VDD pch W=2.8U L=0.24U
M5 Q DIN1 VSS VSS nch W=0.6U L=0.24U
M4 Q DIN1 N1N490 VDD pch W=2.7U L=0.24U
M1 N1N490 DIN2 VDD VDD pch W=2.8U L=0.24U
M3 VDD DIN4 N1N490 VDD pch W=2.8U L=0.24U
M8 VSS DIN4 N1N454 VSS nch W=1U L=0.24U
M7 N1N454 DIN3 N1N452 VSS nch W=1.24U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi13s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 VSS VSS nch W=0.8U L=0.24U
M4 Q DIN1 N1N486 VDD pch W=4U L=0.24U
M1 N1N486 DIN2 VDD VDD pch W=4.1U L=0.24U
M2 VDD DIN3 N1N486 VDD pch W=4.1U L=0.24U
M3 VDD DIN4 N1N486 VDD pch W=4.1U L=0.24U
M6 N1N452 DIN2 Q VSS nch W=1.84U L=0.24U
M7 N1N454 DIN3 N1N452 VSS nch W=1.84U L=0.24U
M8 VSS DIN4 N1N454 VSS nch W=1.84U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi13s3 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 VSS VSS nch W=1U L=0.24U
M4 Q DIN1 N1N486 VDD pch W=6U L=0.24U
M1 N1N486 DIN2 VDD VDD pch W=6U L=0.24U
M2 VDD DIN3 N1N486 VDD pch W=6U L=0.24U
M3 VDD DIN4 N1N486 VDD pch W=6U L=0.24U
M6 N1N452 DIN2 Q VSS nch W=2.8U L=0.24U
M7 N1N454 DIN3 N1N452 VSS nch W=2.8U L=0.24U
M8 VSS DIN4 N1N454 VSS nch W=2.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi211s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N444 VSS nch W=1U L=0.24U
M3 N1N439 DIN4 N1N477 VDD pch W=3.7U L=0.24U
M4 Q DIN3 N1N477 VDD pch W=3.7U L=0.24U
M2 VDD DIN2 N1N439 VDD pch W=3.8U L=0.24U
M1 N1N439 DIN1 VDD VDD pch W=3.8U L=0.24U
M7 Q DIN3 VSS VSS nch W=0.6U L=0.24U
M8 VSS DIN4 Q VSS nch W=0.6U L=0.24U
M6 N1N444 DIN2 VSS VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi211s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N444 VSS nch W=1.3U L=0.24U
M3 N1N439 DIN4 N1N477 VDD pch W=4.8U L=0.24U
M4 Q DIN3 N1N477 VDD pch W=4.7U L=0.24U
M2 VDD DIN2 N1N439 VDD pch W=4.9U L=0.24U
M1 N1N439 DIN1 VDD VDD pch W=4.9U L=0.24U
M7 Q DIN3 VSS VSS nch W=0.8U L=0.24U
M8 VSS DIN4 Q VSS nch W=0.8U L=0.24U
M6 N1N444 DIN2 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi211s3 Q DIN1 DIN2 DIN3 DIN4
M5 N1N467 DIN1 N1N444 VSS nch W=1.4U L=0.24U
M3 N1N439 DIN4 N1N480 VDD pch W=4.1U L=0.24U
M4 N1N467 DIN3 N1N480 VDD pch W=3.9U L=0.24U
M2 VDD DIN2 N1N439 VDD pch W=4.3U L=0.24U
M1 N1N439 DIN1 VDD VDD pch W=4.3U L=0.24U
M7 N1N467 DIN3 VSS VSS nch W=0.7U L=0.24U
M8 VSS DIN4 N1N467 VSS nch W=0.7U L=0.24U
M6 N1N444 DIN2 VSS VSS nch W=1.4U L=0.24U
M9 N1N489 N1N467 VDD VDD pch W=2.4U L=0.24U
M10 N1N489 N1N467 VSS VSS nch W=1.6U L=0.24U
M12 Q N1N489 VSS VSS nch W=2U L=0.24U
M11 Q N1N489 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi21s1 Q DIN1 DIN2 DIN3
M5 Q DIN3 VSS VSS nch W=0.6U L=0.24U
M2 VDD DIN1 N1N344 VDD pch W=2.76U L=0.24U
M3 Q DIN3 N1N344 VDD pch W=2.76U L=0.24U
M1 N1N344 DIN2 VDD VDD pch W=2.76U L=0.24U
M4 Q DIN2 N1N322 VSS nch W=1U L=0.24U
M6 N1N322 DIN1 VSS VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi21s2 Q DIN1 DIN2 DIN3
M5 Q DIN3 VSS VSS nch W=0.8U L=0.24U
M2 VDD DIN1 N1N344 VDD pch W=3.54U L=0.24U
M3 Q DIN3 N1N344 VDD pch W=3.54U L=0.24U
M1 N1N344 DIN2 VDD VDD pch W=3.54U L=0.24U
M4 Q DIN2 N1N322 VSS nch W=1.3U L=0.24U
M6 N1N322 DIN1 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi21s3 Q DIN1 DIN2 DIN3
M5 Q DIN3 VSS VSS nch W=1U L=0.24U
M2 VDD DIN1 N1N344 VDD pch W=4.6U L=0.24U
M3 Q DIN3 N1N344 VDD pch W=4.6U L=0.24U
M1 N1N344 DIN2 VDD VDD pch W=4.6U L=0.24U
M4 Q DIN2 N1N322 VSS nch W=1.7U L=0.24U
M6 N1N322 DIN1 VSS VSS nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi221s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N449 VSS nch W=1U L=0.24U
M1 N1N439 DIN3 VDD VDD pch W=3.6U L=0.24U
M2 VDD DIN4 N1N439 VDD pch W=3.6U L=0.24U
M4 N1N439 DIN2 N1N443 VDD pch W=3.5U L=0.24U
M3 N1N443 DIN1 N1N439 VDD pch W=3.5U L=0.24U
M5 Q DIN5 N1N443 VDD pch W=3.4U L=0.24U
M8 N1N451 DIN3 Q VSS nch W=1U L=0.24U
M10 VSS DIN4 N1N451 VSS nch W=1U L=0.24U
M9 N1N449 DIN2 VSS VSS nch W=1U L=0.24U
M7 Q DIN5 VSS VSS nch W=0.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi221s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N449 VSS nch W=1.22U L=0.24U
M1 N1N439 DIN3 VDD VDD pch W=4.3U L=0.24U
M3 N1N443 DIN1 N1N439 VDD pch W=4.2U L=0.24U
M5 Q DIN5 N1N443 VDD pch W=4.1U L=0.24U
M2 VDD DIN4 N1N439 VDD pch W=4.3U L=0.24U
M4 N1N439 DIN2 N1N443 VDD pch W=4.2U L=0.24U
M9 N1N449 DIN2 VSS VSS nch W=1.22U L=0.24U
M7 Q DIN5 VSS VSS nch W=0.74U L=0.24U
M8 N1N451 DIN3 Q VSS nch W=1.22U L=0.24U
M10 VSS DIN4 N1N451 VSS nch W=1.22U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi221s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N446 DIN1 N1N449 VSS nch W=1.3U L=0.24U
M1 N1N439 DIN3 VDD VDD pch W=3.7U L=0.24U
M3 N1N443 DIN1 N1N439 VDD pch W=3.5U L=0.24U
M5 N1N446 DIN5 N1N443 VDD pch W=3.4U L=0.24U
M2 VDD DIN4 N1N439 VDD pch W=3.7U L=0.24U
M4 N1N439 DIN2 N1N443 VDD pch W=3.5U L=0.24U
M9 N1N449 DIN2 VSS VSS nch W=1.3U L=0.24U
M7 N1N446 DIN5 VSS VSS nch W=0.7U L=0.24U
M8 N1N451 DIN3 N1N446 VSS nch W=1.3U L=0.24U
M10 VSS DIN4 N1N451 VSS nch W=1.3U L=0.24U
M11 N1N527 N1N446 VDD VDD pch W=2.5U L=0.24U
M12 N1N527 N1N446 VSS VSS nch W=1.6U L=0.24U
M14 Q N1N527 VSS VSS nch W=2U L=0.24U
M13 Q N1N527 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi2221s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M1 N1N487 DIN1 VDD VDD pch W=5.8U L=0.24U
M3 N1N489 DIN3 N1N487 VDD pch W=5.6U L=0.24U
M5 N1N452 DIN5 N1N489 VDD pch W=5.4U L=0.24U
M2 VDD DIN2 N1N487 VDD pch W=5.8U L=0.24U
M4 N1N487 DIN4 N1N489 VDD pch W=5.6U L=0.24U
M6 N1N489 DIN6 N1N452 VDD pch W=5.4U L=0.24U
M8 Q DIN1 N1N454 VSS nch W=1.2U L=0.24U
M9 Q DIN3 N1N506 VSS nch W=1.2U L=0.24U
M13 N1N506 DIN4 VSS VSS nch W=1.2U L=0.24U
M12 N1N454 DIN2 VSS VSS nch W=1.2U L=0.24U
M10 N1N508 DIN5 Q VSS nch W=1.2U L=0.24U
M14 VSS DIN6 N1N508 VSS nch W=1.2U L=0.24U
M11 VSS DIN7 Q VSS nch W=0.6U L=0.24U
M7 Q DIN7 N1N452 VDD pch W=5.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi2221s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M1 N1N487 DIN1 VDD VDD pch W=7.1U L=0.24U
M3 N1N489 DIN3 N1N487 VDD pch W=6.9U L=0.24U
M5 N1N452 DIN5 N1N489 VDD pch W=6.7U L=0.24U
M2 VDD DIN2 N1N487 VDD pch W=7.1U L=0.24U
M4 N1N487 DIN4 N1N489 VDD pch W=6.9U L=0.24U
M6 N1N489 DIN6 N1N452 VDD pch W=6.7U L=0.24U
M8 Q DIN1 N1N454 VSS nch W=1.4U L=0.24U
M9 Q DIN3 N1N506 VSS nch W=1.4U L=0.24U
M13 N1N506 DIN4 VSS VSS nch W=1.4U L=0.24U
M12 N1N454 DIN2 VSS VSS nch W=1.4U L=0.24U
M10 N1N508 DIN5 Q VSS nch W=1.4U L=0.24U
M14 VSS DIN6 N1N508 VSS nch W=1.4U L=0.24U
M11 VSS DIN7 Q VSS nch W=0.7U L=0.24U
M7 Q DIN7 N1N452 VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi2221s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M1 N1N487 DIN1 VDD VDD pch W=8.6U L=0.24U
M3 N1N489 DIN3 N1N487 VDD pch W=8.4U L=0.24U
M5 N1N452 DIN5 N1N489 VDD pch W=8.2U L=0.24U
M2 VDD DIN2 N1N487 VDD pch W=8.6U L=0.24U
M4 N1N487 DIN4 N1N489 VDD pch W=8.4U L=0.24U
M6 N1N489 DIN6 N1N452 VDD pch W=8.2U L=0.24U
M8 Q DIN1 N1N454 VSS nch W=1.8U L=0.24U
M9 Q DIN3 N1N506 VSS nch W=1.8U L=0.24U
M13 N1N506 DIN4 VSS VSS nch W=1.8U L=0.24U
M12 N1N454 DIN2 VSS VSS nch W=1.8U L=0.24U
M10 N1N508 DIN5 Q VSS nch W=1.8U L=0.24U
M14 VSS DIN6 N1N508 VSS nch W=1.8U L=0.24U
M11 VSS DIN7 Q VSS nch W=0.9U L=0.24U
M7 Q DIN7 N1N452 VDD pch W=8.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi222s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N453 VSS nch W=1U L=0.24U
M1 N1N441 DIN6 VDD VDD pch W=3.76U L=0.24U
M2 VDD DIN5 N1N441 VDD pch W=3.76U L=0.24U
M3 N1N443 DIN4 N1N441 VDD pch W=3.46U L=0.24U
M4 N1N441 DIN3 N1N443 VDD pch W=3.46U L=0.24U
M5 Q DIN1 N1N443 VDD pch W=3.2U L=0.24U
M6 N1N443 DIN2 Q VDD pch W=3.2U L=0.24U
M10 N1N453 DIN2 VSS VSS nch W=1.1U L=0.24U
M8 Q DIN3 N1N517 VSS nch W=1U L=0.24U
M11 N1N517 DIN4 VSS VSS nch W=1.1U L=0.24U
M9 N1N455 DIN5 Q VSS nch W=1U L=0.24U
M12 VSS DIN6 N1N455 VSS nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi222s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N453 VSS nch W=1.2U L=0.24U
M1 N1N441 DIN6 VDD VDD pch W=4.6U L=0.24U
M2 VDD DIN5 N1N441 VDD pch W=4.6U L=0.24U
M3 N1N443 DIN4 N1N441 VDD pch W=4.2U L=0.24U
M4 N1N441 DIN3 N1N443 VDD pch W=4.2U L=0.24U
M5 Q DIN1 N1N443 VDD pch W=3.8U L=0.24U
M6 N1N443 DIN2 Q VDD pch W=3.8U L=0.24U
M10 N1N453 DIN2 VSS VSS nch W=1.4U L=0.24U
M8 Q DIN3 N1N474 VSS nch W=1.2U L=0.24U
M11 N1N474 DIN4 VSS VSS nch W=1.4U L=0.24U
M9 N1N455 DIN5 Q VSS nch W=1.2U L=0.24U
M12 VSS DIN6 N1N455 VSS nch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi222s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N449 DIN1 N1N453 VSS nch W=1.3U L=0.24U
M1 N1N441 DIN6 VDD VDD pch W=3.8U L=0.24U
M3 N1N443 DIN4 N1N441 VDD pch W=3.6U L=0.24U
M5 N1N449 DIN1 N1N443 VDD pch W=3.3U L=0.24U
M2 VDD DIN5 N1N441 VDD pch W=3.8U L=0.24U
M4 N1N441 DIN3 N1N443 VDD pch W=3.6U L=0.24U
M6 N1N443 DIN2 N1N449 VDD pch W=3.3U L=0.24U
M10 N1N453 DIN2 VSS VSS nch W=1.3U L=0.24U
M8 N1N449 DIN3 N1N474 VSS nch W=1.3U L=0.24U
M11 N1N474 DIN4 VSS VSS nch W=1.3U L=0.24U
M9 N1N455 DIN5 N1N449 VSS nch W=1.3U L=0.24U
M12 VSS DIN6 N1N455 VSS nch W=1.3U L=0.24U
M14 N1N517 N1N449 VSS VSS nch W=1.6U L=0.24U
M13 N1N517 N1N449 VDD VDD pch W=2.8U L=0.24U
M15 Q N1N517 VDD VDD pch W=4.7U L=0.24U
M16 Q N1N517 VSS VSS nch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi22s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N445 VSS nch W=1U L=0.24U
M1 N1N477 DIN3 VDD VDD pch W=2.6U L=0.24U
M3 Q DIN1 N1N477 VDD pch W=2.6U L=0.24U
M2 VDD DIN4 N1N477 VDD pch W=2.6U L=0.24U
M4 N1N477 DIN2 Q VDD pch W=2.6U L=0.24U
M7 N1N445 DIN2 VSS VSS nch W=1U L=0.24U
M6 N1N447 DIN3 Q VSS nch W=1U L=0.24U
M8 VSS DIN4 N1N447 VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi22s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N445 VSS nch W=1.3U L=0.24U
M1 N1N477 DIN3 VDD VDD pch W=3.3U L=0.24U
M3 Q DIN1 N1N477 VDD pch W=3.3U L=0.24U
M2 VDD DIN4 N1N477 VDD pch W=3.3U L=0.24U
M4 N1N477 DIN2 Q VDD pch W=3.3U L=0.24U
M7 N1N445 DIN2 VSS VSS nch W=1.3U L=0.24U
M6 N1N447 DIN3 Q VSS nch W=1.3U L=0.24U
M8 VSS DIN4 N1N447 VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi22s3 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N445 VSS nch W=1.84U L=0.24U
M1 N1N477 DIN3 VDD VDD pch W=4.6U L=0.24U
M3 Q DIN1 N1N477 VDD pch W=4.6U L=0.24U
M2 VDD DIN4 N1N477 VDD pch W=4.6U L=0.24U
M4 N1N477 DIN2 Q VDD pch W=4.6U L=0.24U
M7 N1N445 DIN2 VSS VSS nch W=1.84U L=0.24U
M6 N1N447 DIN3 Q VSS nch W=1.84U L=0.24U
M8 VSS DIN4 N1N447 VSS nch W=1.84U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi23s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N497 VSS nch W=1U L=0.24U
M1 N1N487 DIN3 VDD VDD pch W=2.66U L=0.24U
M3 VDD DIN5 N1N487 VDD pch W=2.66U L=0.24U
M5 N1N487 DIN2 Q VDD pch W=2.6U L=0.24U
M4 Q DIN1 N1N487 VDD pch W=2.6U L=0.24U
M7 N1N497 DIN2 VSS VSS nch W=1U L=0.24U
M10 VSS DIN5 N1N501 VSS nch W=1.3U L=0.24U
M9 N1N501 DIN4 N1N499 VSS nch W=1.3U L=0.24U
M8 N1N499 DIN3 Q VSS nch W=1.3U L=0.24U
M2 VDD DIN4 N1N487 VDD pch W=2.66U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi23s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M2 VDD DIN4 N1N435 VDD pch W=3.5U L=0.24U
M1 N1N435 DIN3 VDD VDD pch W=3.5U L=0.24U
M5 N1N435 DIN2 Q VDD pch W=3.4U L=0.24U
M4 Q DIN1 N1N435 VDD pch W=3.4U L=0.24U
M3 VDD DIN5 N1N435 VDD pch W=3.5U L=0.24U
M6 Q DIN1 N1N463 VSS nch W=1.4U L=0.24U
M7 N1N463 DIN2 VSS VSS nch W=1.4U L=0.24U
M10 VSS DIN5 N1N467 VSS nch W=1.8U L=0.24U
M8 N1N465 DIN3 Q VSS nch W=1.7U L=0.24U
M9 N1N467 DIN4 N1N465 VSS nch W=1.76U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi23s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M2 VDD DIN4 N1N435 VDD pch W=4.8U L=0.24U
M1 N1N435 DIN3 VDD VDD pch W=4.8U L=0.24U
M5 N1N435 DIN2 Q VDD pch W=4.6U L=0.24U
M4 Q DIN1 N1N435 VDD pch W=4.6U L=0.24U
M3 VDD DIN5 N1N435 VDD pch W=4.8U L=0.24U
M6 Q DIN1 N1N463 VSS nch W=1.9U L=0.24U
M7 N1N463 DIN2 VSS VSS nch W=1.9U L=0.24U
M10 VSS DIN5 N1N467 VSS nch W=2.5U L=0.24U
M8 N1N465 DIN3 Q VSS nch W=2.3U L=0.24U
M9 N1N467 DIN4 N1N465 VSS nch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi33s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN6 N1N481 VSS nch W=1.7U L=0.24U
M1 N1N459 DIN2 VDD VDD pch W=2.56U L=0.24U
M4 Q DIN5 N1N459 VDD pch W=2.4U L=0.24U
M2 N1N459 DIN3 VDD VDD pch W=2.56U L=0.24U
M5 Q DIN6 N1N459 VDD pch W=2.4U L=0.24U
M3 VDD DIN1 N1N459 VDD pch W=2.56U L=0.24U
M6 N1N459 DIN4 Q VDD pch W=2.4U L=0.24U
M9 N1N481 DIN5 N1N483 VSS nch W=1.7U L=0.24U
M11 N1N483 DIN4 VSS VSS nch W=1.7U L=0.24U
M10 N1N487 DIN2 N1N485 VSS nch W=1.7U L=0.24U
M8 Q DIN3 N1N485 VSS nch W=1.7U L=0.24U
M12 VSS DIN1 N1N487 VSS nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi33s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN6 N1N481 VSS nch W=2U L=0.24U
M1 N1N459 DIN2 VDD VDD pch W=3.5U L=0.24U
M2 N1N459 DIN3 VDD VDD pch W=3.5U L=0.24U
M4 Q DIN5 N1N459 VDD pch W=3.4U L=0.24U
M5 Q DIN6 N1N459 VDD pch W=3.4U L=0.24U
M3 VDD DIN1 N1N459 VDD pch W=3.5U L=0.24U
M6 N1N459 DIN4 Q VDD pch W=3.4U L=0.24U
M9 N1N481 DIN5 N1N483 VSS nch W=2.5U L=0.24U
M11 N1N483 DIN4 VSS VSS nch W=2.9U L=0.24U
M10 N1N487 DIN2 N1N485 VSS nch W=2.5U L=0.24U
M8 Q DIN3 N1N485 VSS nch W=2U L=0.24U
M12 VSS DIN1 N1N487 VSS nch W=2.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi33s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN6 N1N481 VSS nch W=2.6U L=0.24U
M1 N1N459 DIN2 VDD VDD pch W=4.6U L=0.24U
M4 Q DIN5 N1N459 VDD pch W=4.4U L=0.24U
M2 N1N459 DIN3 VDD VDD pch W=4.6U L=0.24U
M5 Q DIN6 N1N459 VDD pch W=4.4U L=0.24U
M3 VDD DIN1 N1N459 VDD pch W=4.6U L=0.24U
M6 N1N459 DIN4 Q VDD pch W=4.4U L=0.24U
M8 Q DIN3 N1N485 VSS nch W=2.6U L=0.24U
M11 N1N483 DIN4 VSS VSS nch W=3.9U L=0.24U
M10 N1N487 DIN2 N1N485 VSS nch W=3.4U L=0.24U
M9 N1N481 DIN5 N1N483 VSS nch W=3.4U L=0.24U
M12 VSS DIN1 N1N487 VSS nch W=3.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi4111s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 Q DIN7 VSS VSS nch W=0.6U L=0.24U
M5 N1N440 DIN7 N1N613 VDD pch W=5.4U L=0.24U
M6 N1N472 DIN6 N1N440 VDD pch W=5.2U L=0.24U
M7 Q DIN5 N1N472 VDD pch W=5U L=0.24U
M1 N1N613 DIN1 VDD VDD pch W=5.6U L=0.24U
M2 N1N613 DIN2 VDD VDD pch W=5.6U L=0.24U
M3 N1N613 DIN3 VDD VDD pch W=5.6U L=0.24U
M4 N1N613 DIN4 VDD VDD pch W=5.6U L=0.24U
M9 Q DIN6 VSS VSS nch W=0.6U L=0.24U
M10 Q DIN5 VSS VSS nch W=0.6U L=0.24U
M11 Q DIN4 N1N514 VSS nch W=2.4U L=0.24U
M13 N1N515 DIN2 N1N501 VSS nch W=2.4U L=0.24U
M14 N1N501 DIN1 VSS VSS nch W=2.4U L=0.24U
M12 N1N515 DIN3 N1N514 VSS nch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi4111s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 Q DIN7 VSS VSS nch W=0.7U L=0.24U
M5 N1N440 DIN7 N1N613 VDD pch W=6.2U L=0.24U
M6 N1N472 DIN6 N1N440 VDD pch W=6U L=0.24U
M7 Q DIN5 N1N472 VDD pch W=5.8U L=0.24U
M1 N1N613 DIN1 VDD VDD pch W=6.3U L=0.24U
M2 N1N613 DIN2 VDD VDD pch W=6.3U L=0.24U
M3 N1N613 DIN3 VDD VDD pch W=6.3U L=0.24U
M4 N1N613 DIN4 VDD VDD pch W=6.3U L=0.24U
M9 Q DIN6 VSS VSS nch W=0.7U L=0.24U
M10 Q DIN5 VSS VSS nch W=0.7U L=0.24U
M11 Q DIN4 N1N514 VSS nch W=2.8U L=0.24U
M13 N1N515 DIN2 N1N501 VSS nch W=2.8U L=0.24U
M14 N1N501 DIN1 VSS VSS nch W=2.8U L=0.24U
M12 N1N515 DIN3 N1N514 VSS nch W=2.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi4111s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 N1N449 DIN7 VSS VSS nch W=0.6U L=0.24U
M5 N1N440 DIN7 N1N639 VDD pch W=4.8U L=0.24U
M6 N1N472 DIN6 N1N440 VDD pch W=4.6U L=0.24U
M7 N1N449 DIN5 N1N472 VDD pch W=4.4U L=0.24U
M1 N1N639 DIN1 VDD VDD pch W=5U L=0.24U
M2 N1N639 DIN2 VDD VDD pch W=5U L=0.24U
M3 N1N639 DIN3 VDD VDD pch W=5U L=0.24U
M4 N1N639 DIN4 VDD VDD pch W=5U L=0.24U
M9 N1N449 DIN6 VSS VSS nch W=0.6U L=0.24U
M10 N1N449 DIN5 VSS VSS nch W=0.6U L=0.24U
M11 N1N449 DIN4 N1N514 VSS nch W=2.4U L=0.24U
M13 N1N515 DIN2 N1N501 VSS nch W=2.4U L=0.24U
M14 N1N501 DIN1 VSS VSS nch W=2.4U L=0.24U
M12 N1N515 DIN3 N1N514 VSS nch W=2.4U L=0.24U
M16 N1N591 N1N449 VSS VSS nch W=2.2U L=0.24U
M15 N1N591 N1N449 VDD VDD pch W=4.8U L=0.24U
M17 Q N1N591 VDD VDD pch W=6.6U L=0.24U
M18 Q N1N591 VSS VSS nch W=3.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi42s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N447 VSS nch W=1.9U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=2.6U L=0.24U
M2 N1N440 DIN2 VDD VDD pch W=2.6U L=0.24U
M3 VDD DIN3 N1N440 VDD pch W=2.6U L=0.24U
M4 VDD DIN4 N1N440 VDD pch W=2.6U L=0.24U
M5 Q DIN5 N1N440 VDD pch W=2.6U L=0.24U
M6 N1N440 DIN6 Q VDD pch W=2.6U L=0.24U
M8 N1N447 DIN2 N1N463 VSS nch W=1.9U L=0.24U
M9 N1N463 DIN3 N1N465 VSS nch W=1.9U L=0.24U
M10 N1N465 DIN4 VSS VSS nch W=1.9U L=0.24U
M11 N1N451 DIN5 Q VSS nch W=1U L=0.24U
M12 VSS DIN6 N1N451 VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi42s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N447 VSS nch W=2.86U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=3.9U L=0.24U
M2 N1N440 DIN2 VDD VDD pch W=3.9U L=0.24U
M3 VDD DIN3 N1N440 VDD pch W=3.9U L=0.24U
M4 VDD DIN4 N1N440 VDD pch W=3.9U L=0.24U
M5 Q DIN5 N1N440 VDD pch W=3.9U L=0.24U
M6 N1N440 DIN6 Q VDD pch W=3.9U L=0.24U
M8 N1N447 DIN2 N1N463 VSS nch W=2.86U L=0.24U
M9 N1N463 DIN3 N1N465 VSS nch W=2.86U L=0.24U
M10 N1N465 DIN4 VSS VSS nch W=2.86U L=0.24U
M11 N1N451 DIN5 Q VSS nch W=1.5U L=0.24U
M12 VSS DIN6 N1N451 VSS nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT aoi42s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N447 VSS nch W=4.3U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=5.9U L=0.24U
M2 N1N440 DIN2 VDD VDD pch W=5.9U L=0.24U
M3 VDD DIN3 N1N440 VDD pch W=5.9U L=0.24U
M4 VDD DIN4 N1N440 VDD pch W=5.9U L=0.24U
M5 Q DIN5 N1N440 VDD pch W=5.9U L=0.24U
M6 N1N440 DIN6 Q VDD pch W=5.9U L=0.24U
M8 N1N447 DIN2 N1N463 VSS nch W=4.3U L=0.24U
M9 N1N463 DIN3 N1N465 VSS nch W=4.3U L=0.24U
M10 N1N465 DIN4 VSS VSS nch W=4.3U L=0.24U
M11 N1N451 DIN5 Q VSS nch W=2.26U L=0.24U
M12 VSS DIN6 N1N451 VSS nch W=2.26U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT bshes1 INOUT1 INOUT2 E
M2 N1N313 E VSS VSS nch W=0.8U L=0.24U
M1 N1N313 E VDD VDD pch W=1.2U L=0.24U
M3 INOUT2 N1N313 INOUT1 VDD pch W=1.2U L=0.24U
M4 INOUT1 E INOUT2 VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT bshes2 INOUT2 E INOUT1
M2 N1N313 E VSS VSS nch W=1U L=0.24U
M1 N1N313 E VDD VDD pch W=1.5U L=0.24U
M3 INOUT2 N1N313 INOUT1 VDD pch W=2.1U L=0.24U
M4 INOUT1 E INOUT2 VSS nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT bshes3 INOUT2 E INOUT1
M2 N1N313 E VSS VSS nch W=1.2U L=0.24U
M1 N1N313 E VDD VDD pch W=2U L=0.24U
M3 INOUT2 N1N313 INOUT1 VDD pch W=3.5U L=0.24U
M4 INOUT1 E INOUT2 VSS nch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT bsles1 INOUT2 EB INOUT1
M2 N1N330 EB VSS VSS nch W=0.9U L=0.24U
M1 N1N330 EB VDD VDD pch W=1.15U L=0.24U
M3 INOUT2 EB INOUT1 VDD pch W=1.45U L=0.24U
M4 INOUT1 N1N330 INOUT2 VSS nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT bsles2 INOUT2 EB INOUT1
M2 N1N330 EB VSS VSS nch W=1U L=0.24U
M1 N1N330 EB VDD VDD pch W=1.5U L=0.24U
M3 INOUT2 EB INOUT1 VDD pch W=2.1U L=0.24U
M4 INOUT1 N1N330 INOUT2 VSS nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT bsles3 INOUT2 EB INOUT1
M2 N1N330 EB VSS VSS nch W=1.2U L=0.24U
M1 N1N330 EB VDD VDD pch W=2U L=0.24U
M3 INOUT2 EB INOUT1 VDD pch W=3.5U L=0.24U
M4 INOUT1 N1N330 INOUT2 VSS nch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT clc2s1 PIN0 CIN0 GIN0 GIN1 PIN1 OUTP OUTC OUTG
M14 OUTC N1N64 VSS VSS nch W=0.72U L=0.24U
M7 OUTC N1N64 VDD VDD pch W=1.4U L=0.24U
M16 OUTG N1N145 VSS VSS nch W=0.72U L=0.24U
M15 OUTG N1N145 VDD VDD pch W=1.4U L=0.24U
M17 N1N153 PIN0 VDD VDD pch W=0.9U L=0.24U
M18 N1N153 PIN1 VDD VDD pch W=0.9U L=0.24U
M19 N1N153 PIN0 N1N151 VSS nch W=0.7U L=0.24U
M20 N1N151 PIN1 VSS VSS nch W=0.7U L=0.24U
M22 OUTP N1N153 VSS VSS nch W=0.9U L=0.24U
M21 OUTP N1N153 VDD VDD pch W=1.76U L=0.24U
M6 VSS PIN0 N1N66 VSS nch W=1.2U L=0.24U
M4 N1N64 GIN0 VSS VSS nch W=0.6U L=0.24U
M5 N1N66 CIN0 N1N64 VSS nch W=1.2U L=0.24U
M1 N1N60 PIN0 VDD VDD pch W=2.7U L=0.24U
M2 VDD CIN0 N1N60 VDD pch W=2.7U L=0.24U
M3 N1N64 GIN0 N1N60 VDD pch W=2.7U L=0.24U
M8 N1N86 GIN0 VDD VDD pch W=2.7U L=0.24U
M9 VDD PIN1 N1N86 VDD pch W=2.7U L=0.24U
M10 N1N145 GIN1 N1N86 VDD pch W=2.7U L=0.24U
M11 N1N145 GIN1 VSS VSS nch W=0.6U L=0.24U
M12 N1N85 PIN1 N1N145 VSS nch W=1.2U L=0.24U
M13 VSS GIN0 N1N85 VSS nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT clc2s2 PIN0 CIN0 GIN0 GIN1 PIN1 OUTP OUTC OUTG
M14 OUTC N1N64 VSS VSS nch W=0.92U L=0.24U
M7 OUTC N1N64 VDD VDD pch W=1.7U L=0.24U
M16 OUTG N1N145 VSS VSS nch W=0.92U L=0.24U
M15 OUTG N1N145 VDD VDD pch W=1.7U L=0.24U
M17 N1N153 PIN0 VDD VDD pch W=1.2U L=0.24U
M18 N1N153 PIN1 VDD VDD pch W=1.2U L=0.24U
M19 N1N153 PIN0 N1N151 VSS nch W=0.9U L=0.24U
M20 N1N151 PIN1 VSS VSS nch W=0.9U L=0.24U
M22 OUTP N1N153 VSS VSS nch W=1.2U L=0.24U
M21 OUTP N1N153 VDD VDD pch W=2.26U L=0.24U
M6 VSS PIN0 N1N66 VSS nch W=1.6U L=0.24U
M4 N1N64 GIN0 VSS VSS nch W=0.8U L=0.24U
M5 N1N66 CIN0 N1N64 VSS nch W=1.6U L=0.24U
M1 N1N60 PIN0 VDD VDD pch W=3.5U L=0.24U
M2 VDD CIN0 N1N60 VDD pch W=3.5U L=0.24U
M3 N1N64 GIN0 N1N60 VDD pch W=3.5U L=0.24U
M8 N1N86 GIN0 VDD VDD pch W=3.5U L=0.24U
M9 VDD PIN1 N1N86 VDD pch W=3.5U L=0.24U
M10 N1N145 GIN1 N1N86 VDD pch W=3.5U L=0.24U
M11 N1N145 GIN1 VSS VSS nch W=0.8U L=0.24U
M12 N1N85 PIN1 N1N145 VSS nch W=1.6U L=0.24U
M13 VSS GIN0 N1N85 VSS nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT clc2s3 PIN0 CIN0 GIN0 GIN1 PIN1 OUTP OUTC OUTG
M14 OUTC N1N64 VSS VSS nch W=1.26U L=0.24U
M7 OUTC N1N64 VDD VDD pch W=2.2U L=0.24U
M16 OUTG N1N145 VSS VSS nch W=1.26U L=0.24U
M15 OUTG N1N145 VDD VDD pch W=2.2U L=0.24U
M17 N1N153 PIN0 VDD VDD pch W=1.74U L=0.24U
M18 N1N153 PIN1 VDD VDD pch W=1.74U L=0.24U
M19 N1N153 PIN0 N1N151 VSS nch W=1.2U L=0.24U
M20 N1N151 PIN1 VSS VSS nch W=1.2U L=0.24U
M22 OUTP N1N153 VSS VSS nch W=1.5U L=0.24U
M21 OUTP N1N153 VDD VDD pch W=2.9U L=0.24U
M6 VSS PIN0 N1N66 VSS nch W=2U L=0.24U
M4 N1N64 GIN0 VSS VSS nch W=1U L=0.24U
M5 N1N66 CIN0 N1N64 VSS nch W=2U L=0.24U
M1 N1N60 PIN0 VDD VDD pch W=4.9U L=0.24U
M2 VDD CIN0 N1N60 VDD pch W=4.9U L=0.24U
M3 N1N64 GIN0 N1N60 VDD pch W=4.7U L=0.24U
M8 N1N86 GIN0 VDD VDD pch W=4.9U L=0.24U
M9 VDD PIN1 N1N86 VDD pch W=4.9U L=0.24U
M10 N1N145 GIN1 N1N86 VDD pch W=4.7U L=0.24U
M11 N1N145 GIN1 VSS VSS nch W=1U L=0.24U
M12 N1N85 PIN1 N1N145 VSS nch W=2U L=0.24U
M13 VSS GIN0 N1N85 VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dchei24s1 BIN0 BIN1 E OUTD0 OUTD1 OUTD2 OUTD3
M15 OUTD1 N1N430 VDD VDD pch W=1.3U L=0.24U
M17 OUTD1 N1N301 VDD VDD pch W=1.3U L=0.24U
M20 N1N293 N1N301 VSS VSS nch W=1.16U L=0.24U
M19 N1N294 BIN0 N1N293 VSS nch W=1.16U L=0.24U
M18 OUTD1 N1N430 N1N294 VSS nch W=1.16U L=0.24U
M16 OUTD1 BIN0 VDD VDD pch W=1.3U L=0.24U
M21 OUTD2 N1N430 VDD VDD pch W=1.3U L=0.24U
M23 OUTD2 BIN1 VDD VDD pch W=1.3U L=0.24U
M26 N1N325 BIN1 VSS VSS nch W=1.16U L=0.24U
M25 N1N324 N1N290 N1N325 VSS nch W=1.16U L=0.24U
M24 OUTD2 N1N430 N1N324 VSS nch W=1.16U L=0.24U
M22 OUTD2 N1N290 VDD VDD pch W=1.3U L=0.24U
M9 OUTD0 N1N430 VDD VDD pch W=1.3U L=0.24U
M11 OUTD0 N1N301 VDD VDD pch W=1.3U L=0.24U
M14 N1N344 N1N301 VSS VSS nch W=1.16U L=0.24U
M13 N1N343 N1N290 N1N344 VSS nch W=1.16U L=0.24U
M12 OUTD0 N1N430 N1N343 VSS nch W=1.16U L=0.24U
M10 OUTD0 N1N290 VDD VDD pch W=1.3U L=0.24U
M27 OUTD3 N1N430 VDD VDD pch W=1.3U L=0.24U
M29 OUTD3 BIN1 VDD VDD pch W=1.3U L=0.24U
M32 N1N363 BIN1 VSS VSS nch W=1.16U L=0.24U
M31 N1N362 BIN0 N1N363 VSS nch W=1.16U L=0.24U
M30 OUTD3 N1N430 N1N362 VSS nch W=1.16U L=0.24U
M28 OUTD3 BIN0 VDD VDD pch W=1.3U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M2 N1N301 BIN1 VSS VSS nch W=0.9U L=0.24U
M3 N1N290 BIN0 VDD VDD pch W=1.8U L=0.24U
M4 N1N290 BIN0 VSS VSS nch W=0.9U L=0.24U
M5 N1N384 E VDD VDD pch W=1.2U L=0.24U
M7 N1N430 N1N384 VDD VDD pch W=1.6U L=0.24U
M6 N1N384 E VSS VSS nch W=0.6U L=0.24U
M8 N1N430 N1N384 VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dchei24s2 BIN0 BIN1 E OUTD0 OUTD1 OUTD2 OUTD3
M15 OUTD1 N1N430 VDD VDD pch W=2U L=0.24U
M17 OUTD1 N1N301 VDD VDD pch W=2U L=0.24U
M20 N1N293 N1N301 VSS VSS nch W=1.86U L=0.24U
M19 N1N294 BIN0 N1N293 VSS nch W=1.86U L=0.24U
M18 OUTD1 N1N430 N1N294 VSS nch W=1.86U L=0.24U
M16 OUTD1 BIN0 VDD VDD pch W=2U L=0.24U
M21 OUTD2 N1N430 VDD VDD pch W=2U L=0.24U
M23 OUTD2 BIN1 VDD VDD pch W=2U L=0.24U
M26 N1N325 BIN1 VSS VSS nch W=1.86U L=0.24U
M25 N1N324 N1N290 N1N325 VSS nch W=1.86U L=0.24U
M24 OUTD2 N1N430 N1N324 VSS nch W=1.86U L=0.24U
M22 OUTD2 N1N290 VDD VDD pch W=2U L=0.24U
M9 OUTD0 N1N430 VDD VDD pch W=2U L=0.24U
M11 OUTD0 N1N301 VDD VDD pch W=2U L=0.24U
M14 N1N344 N1N301 VSS VSS nch W=1.86U L=0.24U
M13 N1N343 N1N290 N1N344 VSS nch W=1.86U L=0.24U
M12 OUTD0 N1N430 N1N343 VSS nch W=1.86U L=0.24U
M10 OUTD0 N1N290 VDD VDD pch W=2U L=0.24U
M27 OUTD3 N1N430 VDD VDD pch W=2U L=0.24U
M29 OUTD3 BIN1 VDD VDD pch W=2U L=0.24U
M32 N1N363 BIN1 VSS VSS nch W=1.86U L=0.24U
M31 N1N362 BIN0 N1N363 VSS nch W=1.86U L=0.24U
M30 OUTD3 N1N430 N1N362 VSS nch W=1.86U L=0.24U
M28 OUTD3 BIN0 VDD VDD pch W=2U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M2 N1N301 BIN1 VSS VSS nch W=0.8U L=0.24U
M3 N1N290 BIN0 VDD VDD pch W=1.8U L=0.24U
M4 N1N290 BIN0 VSS VSS nch W=0.9U L=0.24U
M5 N1N384 E VDD VDD pch W=1.2U L=0.24U
M7 N1N430 N1N384 VDD VDD pch W=1.6U L=0.24U
M6 N1N384 E VSS VSS nch W=0.6U L=0.24U
M8 N1N430 N1N384 VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dchei24s3 BIN0 BIN1 E OUTD0 OUTD1 OUTD2 OUTD3
M15 OUTD1 N1N430 VDD VDD pch W=3U L=0.24U
M17 OUTD1 N1N301 VDD VDD pch W=3U L=0.24U
M20 N1N293 N1N301 VSS VSS nch W=2.92U L=0.24U
M19 N1N294 BIN0 N1N293 VSS nch W=2.92U L=0.24U
M18 OUTD1 N1N430 N1N294 VSS nch W=2.92U L=0.24U
M16 OUTD1 BIN0 VDD VDD pch W=3U L=0.24U
M21 OUTD2 N1N430 VDD VDD pch W=3U L=0.24U
M23 OUTD2 BIN1 VDD VDD pch W=3U L=0.24U
M26 N1N325 BIN1 VSS VSS nch W=2.92U L=0.24U
M25 N1N324 N1N290 N1N325 VSS nch W=2.92U L=0.24U
M24 OUTD2 N1N430 N1N324 VSS nch W=2.92U L=0.24U
M22 OUTD2 N1N290 VDD VDD pch W=3U L=0.24U
M9 OUTD0 N1N430 VDD VDD pch W=3U L=0.24U
M11 OUTD0 N1N301 VDD VDD pch W=3U L=0.24U
M14 N1N344 N1N301 VSS VSS nch W=2.92U L=0.24U
M13 N1N343 N1N290 N1N344 VSS nch W=2.92U L=0.24U
M12 OUTD0 N1N430 N1N343 VSS nch W=2.92U L=0.24U
M10 OUTD0 N1N290 VDD VDD pch W=3U L=0.24U
M27 OUTD3 N1N430 VDD VDD pch W=3U L=0.24U
M29 OUTD3 BIN1 VDD VDD pch W=3U L=0.24U
M32 N1N363 BIN1 VSS VSS nch W=2.92U L=0.24U
M31 N1N362 BIN0 N1N363 VSS nch W=2.92U L=0.24U
M30 OUTD3 N1N430 N1N362 VSS nch W=2.92U L=0.24U
M28 OUTD3 BIN0 VDD VDD pch W=3U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M2 N1N301 BIN1 VSS VSS nch W=0.8U L=0.24U
M3 N1N290 BIN0 VDD VDD pch W=1.8U L=0.24U
M4 N1N290 BIN0 VSS VSS nch W=0.9U L=0.24U
M5 N1N384 E VDD VDD pch W=1.2U L=0.24U
M7 N1N430 N1N384 VDD VDD pch W=1.6U L=0.24U
M6 N1N384 E VSS VSS nch W=0.6U L=0.24U
M8 N1N430 N1N384 VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dci24s1 OUTD0 OUTD1 OUTD2 OUTD3 BIN1 BIN0
M2 N1N301 BIN1 VSS VSS nch W=0.9U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N404 BIN0 VSS VSS nch W=0.9U L=0.24U
M3 N1N404 BIN0 VDD VDD pch W=1.8U L=0.24U
M5 OUTD0 N1N404 VDD VDD pch W=1.66U L=0.24U
M6 VDD N1N301 OUTD0 VDD pch W=1.66U L=0.24U
M7 OUTD0 N1N404 N1N344 VSS nch W=1.2U L=0.24U
M8 N1N344 N1N301 VSS VSS nch W=1.2U L=0.24U
M12 N1N341 N1N301 VSS VSS nch W=1.2U L=0.24U
M11 OUTD1 BIN0 N1N341 VSS nch W=1.2U L=0.24U
M10 VDD N1N301 OUTD1 VDD pch W=1.66U L=0.24U
M9 OUTD1 BIN0 VDD VDD pch W=1.66U L=0.24U
M16 N1N338 N1N404 VSS VSS nch W=1.2U L=0.24U
M15 OUTD2 BIN1 N1N338 VSS nch W=1.2U L=0.24U
M14 VDD N1N404 OUTD2 VDD pch W=1.66U L=0.24U
M13 OUTD2 BIN1 VDD VDD pch W=1.66U L=0.24U
M20 N1N335 BIN1 VSS VSS nch W=1.2U L=0.24U
M19 OUTD3 BIN0 N1N335 VSS nch W=1.2U L=0.24U
M18 VDD BIN1 OUTD3 VDD pch W=1.66U L=0.24U
M17 OUTD3 BIN0 VDD VDD pch W=1.66U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dci24s2 OUTD0 OUTD1 OUTD2 OUTD3 BIN1 BIN0
M2 N1N301 BIN1 VSS VSS nch W=0.9U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N404 BIN0 VSS VSS nch W=0.9U L=0.24U
M3 N1N404 BIN0 VDD VDD pch W=1.8U L=0.24U
M5 OUTD0 N1N404 VDD VDD pch W=2.3U L=0.24U
M6 VDD N1N301 OUTD0 VDD pch W=2.3U L=0.24U
M7 OUTD0 N1N404 N1N344 VSS nch W=1.8U L=0.24U
M8 N1N344 N1N301 VSS VSS nch W=1.8U L=0.24U
M12 N1N341 N1N301 VSS VSS nch W=1.8U L=0.24U
M11 OUTD1 BIN0 N1N341 VSS nch W=1.8U L=0.24U
M10 VDD N1N301 OUTD1 VDD pch W=2.3U L=0.24U
M9 OUTD1 BIN0 VDD VDD pch W=2.3U L=0.24U
M16 N1N338 N1N404 VSS VSS nch W=1.8U L=0.24U
M15 OUTD2 BIN1 N1N338 VSS nch W=1.8U L=0.24U
M14 VDD N1N404 OUTD2 VDD pch W=2.3U L=0.24U
M13 OUTD2 BIN1 VDD VDD pch W=2.3U L=0.24U
M20 N1N335 BIN1 VSS VSS nch W=1.8U L=0.24U
M19 OUTD3 BIN0 N1N335 VSS nch W=1.8U L=0.24U
M18 VDD BIN1 OUTD3 VDD pch W=2.3U L=0.24U
M17 OUTD3 BIN0 VDD VDD pch W=2.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dci24s3 OUTD0 OUTD1 OUTD2 OUTD3 BIN1 BIN0
M2 N1N301 BIN1 VSS VSS nch W=0.9U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N404 BIN0 VSS VSS nch W=0.9U L=0.24U
M3 N1N404 BIN0 VDD VDD pch W=1.8U L=0.24U
M5 OUTD0 N1N404 VDD VDD pch W=4.2U L=0.24U
M6 VDD N1N301 OUTD0 VDD pch W=4.2U L=0.24U
M7 OUTD0 N1N404 N1N344 VSS nch W=4U L=0.24U
M8 N1N344 N1N301 VSS VSS nch W=4U L=0.24U
M12 N1N341 N1N301 VSS VSS nch W=4U L=0.24U
M11 OUTD1 BIN0 N1N341 VSS nch W=4U L=0.24U
M10 VDD N1N301 OUTD1 VDD pch W=4.2U L=0.24U
M9 OUTD1 BIN0 VDD VDD pch W=4.2U L=0.24U
M16 N1N338 N1N404 VSS VSS nch W=4U L=0.24U
M15 OUTD2 BIN1 N1N338 VSS nch W=4U L=0.24U
M14 VDD N1N404 OUTD2 VDD pch W=4.2U L=0.24U
M13 OUTD2 BIN1 VDD VDD pch W=4.2U L=0.24U
M20 N1N335 BIN1 VSS VSS nch W=4U L=0.24U
M19 OUTD3 BIN0 N1N335 VSS nch W=4U L=0.24U
M18 VDD BIN1 OUTD3 VDD pch W=4.2U L=0.24U
M17 OUTD3 BIN0 VDD VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dclei24s1 BIN0 BIN1 EB OUTD0 OUTD1 OUTD2 OUTD3
M10 OUTD0 N1N344 N1N340 VSS nch W=1.16U L=0.24U
M7 OUTD0 N1N344 VDD VDD pch W=1.3U L=0.24U
M8 OUTD0 N1N334 VDD VDD pch W=1.3U L=0.24U
M9 OUTD0 N1N346 VDD VDD pch W=1.3U L=0.24U
M11 N1N340 N1N334 N1N342 VSS nch W=1.16U L=0.24U
M12 N1N342 N1N346 VSS VSS nch W=1.16U L=0.24U
M16 OUTD1 N1N344 N1N373 VSS nch W=1.16U L=0.24U
M13 OUTD1 N1N344 VDD VDD pch W=1.3U L=0.24U
M15 OUTD1 N1N346 VDD VDD pch W=1.3U L=0.24U
M14 OUTD1 BIN0 VDD VDD pch W=1.3U L=0.24U
M17 N1N373 BIN0 N1N374 VSS nch W=1.16U L=0.24U
M18 N1N374 N1N346 VSS VSS nch W=1.16U L=0.24U
M22 OUTD2 N1N344 N1N389 VSS nch W=1.16U L=0.24U
M19 OUTD2 N1N344 VDD VDD pch W=1.3U L=0.24U
M21 OUTD2 BIN1 VDD VDD pch W=1.3U L=0.24U
M20 OUTD2 N1N334 VDD VDD pch W=1.3U L=0.24U
M23 N1N389 N1N334 N1N451 VSS nch W=1.16U L=0.24U
M24 N1N451 BIN1 VSS VSS nch W=1.16U L=0.24U
M28 OUTD3 N1N344 N1N405 VSS nch W=1.16U L=0.24U
M25 OUTD3 N1N344 VDD VDD pch W=1.3U L=0.24U
M27 OUTD3 BIN1 VDD VDD pch W=1.3U L=0.24U
M26 OUTD3 BIN0 VDD VDD pch W=1.3U L=0.24U
M29 N1N405 BIN0 N1N406 VSS nch W=1.16U L=0.24U
M30 N1N406 BIN1 VSS VSS nch W=1.16U L=0.24U
M3 N1N346 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N346 BIN1 VSS VSS nch W=0.9U L=0.24U
M1 N1N334 BIN0 VDD VDD pch W=1.8U L=0.24U
M2 N1N334 BIN0 VSS VSS nch W=0.9U L=0.24U
M6 N1N344 EB VSS VSS nch W=1.2U L=0.24U
M5 N1N344 EB VDD VDD pch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dclei24s2 BIN0 BIN1 EB OUTD0 OUTD1 OUTD2 OUTD3
M10 OUTD0 N1N344 N1N340 VSS nch W=1.86U L=0.24U
M7 OUTD0 N1N344 VDD VDD pch W=2U L=0.24U
M8 OUTD0 N1N334 VDD VDD pch W=2U L=0.24U
M9 OUTD0 N1N346 VDD VDD pch W=2U L=0.24U
M11 N1N340 N1N334 N1N342 VSS nch W=1.86U L=0.24U
M12 N1N342 N1N346 VSS VSS nch W=1.86U L=0.24U
M16 OUTD1 N1N344 N1N373 VSS nch W=1.86U L=0.24U
M13 OUTD1 N1N344 VDD VDD pch W=2U L=0.24U
M15 OUTD1 N1N346 VDD VDD pch W=2U L=0.24U
M14 OUTD1 BIN0 VDD VDD pch W=2U L=0.24U
M17 N1N373 BIN0 N1N374 VSS nch W=1.86U L=0.24U
M18 N1N374 N1N346 VSS VSS nch W=1.86U L=0.24U
M22 OUTD2 N1N344 N1N389 VSS nch W=1.86U L=0.24U
M19 OUTD2 N1N344 VDD VDD pch W=2U L=0.24U
M21 OUTD2 BIN1 VDD VDD pch W=2U L=0.24U
M20 OUTD2 N1N334 VDD VDD pch W=2U L=0.24U
M23 N1N389 N1N334 N1N451 VSS nch W=1.86U L=0.24U
M24 N1N451 BIN1 VSS VSS nch W=1.86U L=0.24U
M28 OUTD3 N1N344 N1N405 VSS nch W=1.86U L=0.24U
M25 OUTD3 N1N344 VDD VDD pch W=2U L=0.24U
M27 OUTD3 BIN1 VDD VDD pch W=2U L=0.24U
M26 OUTD3 BIN0 VDD VDD pch W=2U L=0.24U
M29 N1N405 BIN0 N1N406 VSS nch W=1.86U L=0.24U
M30 N1N406 BIN1 VSS VSS nch W=1.86U L=0.24U
M3 N1N346 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N346 BIN1 VSS VSS nch W=0.9U L=0.24U
M1 N1N334 BIN0 VDD VDD pch W=1.8U L=0.24U
M2 N1N334 BIN0 VSS VSS nch W=0.9U L=0.24U
M6 N1N344 EB VSS VSS nch W=1.2U L=0.24U
M5 N1N344 EB VDD VDD pch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dclei24s3 BIN0 BIN1 EB OUTD0 OUTD1 OUTD2 OUTD3
M10 OUTD0 N1N344 N1N340 VSS nch W=2.94U L=0.24U
M7 OUTD0 N1N344 VDD VDD pch W=3U L=0.24U
M8 OUTD0 N1N334 VDD VDD pch W=3U L=0.24U
M9 OUTD0 N1N346 VDD VDD pch W=3U L=0.24U
M11 N1N340 N1N334 N1N342 VSS nch W=2.94U L=0.24U
M12 N1N342 N1N346 VSS VSS nch W=2.94U L=0.24U
M16 OUTD1 N1N344 N1N373 VSS nch W=2.94U L=0.24U
M13 OUTD1 N1N344 VDD VDD pch W=3U L=0.24U
M15 OUTD1 N1N346 VDD VDD pch W=3U L=0.24U
M14 OUTD1 BIN0 VDD VDD pch W=3U L=0.24U
M17 N1N373 BIN0 N1N374 VSS nch W=2.94U L=0.24U
M18 N1N374 N1N346 VSS VSS nch W=2.94U L=0.24U
M22 OUTD2 N1N344 N1N389 VSS nch W=2.94U L=0.24U
M19 OUTD2 N1N344 VDD VDD pch W=3U L=0.24U
M21 OUTD2 BIN1 VDD VDD pch W=3U L=0.24U
M20 OUTD2 N1N334 VDD VDD pch W=3U L=0.24U
M23 N1N389 N1N334 N1N451 VSS nch W=2.94U L=0.24U
M24 N1N451 BIN1 VSS VSS nch W=2.94U L=0.24U
M28 OUTD3 N1N344 N1N405 VSS nch W=2.94U L=0.24U
M25 OUTD3 N1N344 VDD VDD pch W=3U L=0.24U
M27 OUTD3 BIN1 VDD VDD pch W=3U L=0.24U
M26 OUTD3 BIN0 VDD VDD pch W=3U L=0.24U
M29 N1N405 BIN0 N1N406 VSS nch W=2.94U L=0.24U
M30 N1N406 BIN1 VSS VSS nch W=2.94U L=0.24U
M3 N1N346 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N346 BIN1 VSS VSS nch W=0.9U L=0.24U
M1 N1N334 BIN0 VDD VDD pch W=1.8U L=0.24U
M2 N1N334 BIN0 VSS VSS nch W=0.9U L=0.24U
M6 N1N344 EB VSS VSS nch W=1.2U L=0.24U
M5 N1N344 EB VDD VDD pch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffacs1 Q QN CLRB CLK DIN
M17 TP7 CLRB VDD VDD pch W=1.3U L=0.24U
M21 Q TP8 VDD VDD pch W=3.14U L=0.24U
M9 TP5 TP3 VDD VDD pch W=1.3U L=0.24U
M24 QN Q VSS VSS nch W=1.42U L=0.24U
M3 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M4 DIN TP1 TP3 VSS nch W=0.8U L=0.24U
M13 TP5 CLK TP8 VSS nch W=0.96U L=0.24U
M14 TP8 TP1 TP5 VDD pch W=1.4U L=0.24U
M6 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M15 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M16 TP8 TP1 TP7 VSS nch W=0.8U L=0.24U
M23 QN Q VDD VDD pch W=3.02U L=0.24U
M5 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M11 TP5 TP3 TP6 VSS nch W=0.9U L=0.24U
M19 TP7 Q TP9 VSS nch W=0.9U L=0.24U
M22 Q TP8 VSS VSS nch W=1.96U L=0.24U
M10 TP5 CLRB VDD VDD pch W=1.3U L=0.24U
M8 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M12 TP6 CLRB VSS VSS nch W=0.9U L=0.24U
M1 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M7 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M18 TP7 Q VDD VDD pch W=1.3U L=0.24U
M20 TP9 CLRB VSS VSS nch W=0.9U L=0.24U
M2 TP1 CLK VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffacs2 Q QN CLRB CLK DIN
M17 TP7 CLRB VDD VDD pch W=1.3U L=0.24U
M21 Q TP8 VDD VDD pch W=6.2U L=0.24U
M9 TP5 TP3 VDD VDD pch W=1.84U L=0.24U
M24 QN Q VSS VSS nch W=2.68U L=0.24U
M3 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M4 DIN TP1 TP3 VSS nch W=0.8U L=0.24U
M13 TP5 CLK TP8 VSS nch W=1.52U L=0.24U
M14 TP8 TP1 TP5 VDD pch W=1.9U L=0.24U
M6 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M15 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M16 TP8 TP1 TP7 VSS nch W=0.8U L=0.24U
M23 QN Q VDD VDD pch W=6.16U L=0.24U
M5 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M11 TP5 TP3 TP6 VSS nch W=1.48U L=0.24U
M19 TP7 Q TP9 VSS nch W=0.9U L=0.24U
M22 Q TP8 VSS VSS nch W=3.98U L=0.24U
M10 TP5 CLRB VDD VDD pch W=1.84U L=0.24U
M8 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M12 TP6 CLRB VSS VSS nch W=1.48U L=0.24U
M1 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M7 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M18 TP7 Q VDD VDD pch W=1.3U L=0.24U
M20 TP9 CLRB VSS VSS nch W=0.9U L=0.24U
M2 TP1 CLK VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffascs1 SETB CLRB DIN CLK QN Q
M4 TP2 TP4 VDD VDD pch W=1.8U L=0.24U
M12 TP6 CLK VSS VSS nch W=0.8U L=0.24U
M3 TP2 TP0 VDD VDD pch W=1.8U L=0.24U
M2 TP0 SETB VSS VSS nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M8 TP1 CLRB VSS VSS nch W=0.8U L=0.24U
M7 TP1 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP1 VDD VDD pch W=2.2U L=0.24U
M10 TP4 TP1 VSS VSS nch W=1.4U L=0.24U
M38 QN Q VSS VSS nch W=1.44U L=0.24U
M30 TP14 Q VDD VDD pch W=1.3U L=0.24U
M33 Q TP13 VDD VDD pch W=3.18U L=0.24U
M23 TP11 TP8 TP12 VSS nch W=2.2U L=0.24U
M13 TP8 CLK DIN VDD pch W=1.3U L=0.24U
M14 DIN TP6 TP8 VSS nch W=0.8U L=0.24U
M25 TP11 CLK TP13 VSS nch W=2.2U L=0.24U
M26 TP13 TP6 TP11 VDD pch W=2.5U L=0.24U
M15 TP8 CLK TP9 VSS nch W=0.8U L=0.24U
M16 TP9 TP6 TP8 VDD pch W=1.3U L=0.24U
M27 TP14 CLK TP13 VDD pch W=1.3U L=0.24U
M28 TP13 TP6 TP14 VSS nch W=0.8U L=0.24U
M17 TP9 TP2 VDD VDD pch W=1.3U L=0.24U
M21 TP11 TP8 VDD VDD pch W=2.4U L=0.24U
M22 TP11 TP4 VDD VDD pch W=2.4U L=0.24U
M29 TP14 TP4 VDD VDD pch W=1.3U L=0.24U
M37 QN Q VDD VDD pch W=3.18U L=0.24U
M31 TP14 Q TP15 VSS nch W=0.8U L=0.24U
M20 TP10 TP11 VSS VSS nch W=0.8U L=0.24U
M32 TP15 TP4 VSS VSS nch W=0.8U L=0.24U
M24 TP12 TP4 VSS VSS nch W=2.2U L=0.24U
M36 TP16 TP13 VSS VSS nch W=2.64U L=0.24U
M34 Q TP2 VDD VDD pch W=3.18U L=0.24U
M35 Q TP2 TP16 VSS nch W=2.64U L=0.24U
M18 TP9 TP11 VDD VDD pch W=1.3U L=0.24U
M19 TP9 TP2 TP10 VSS nch W=0.8U L=0.24U
M11 TP6 CLK VDD VDD pch W=1.4U L=0.24U
M5 TP2 TP0 TP3 VSS nch W=1.3U L=0.24U
M6 TP3 TP4 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffascs2 SETB CLRB DIN CLK QN Q
M4 TP2 TP4 VDD VDD pch W=2.82U L=0.24U
M12 TP6 CLK VSS VSS nch W=0.8U L=0.24U
M3 TP2 TP0 VDD VDD pch W=2.82U L=0.24U
M2 TP0 SETB VSS VSS nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M8 TP1 CLRB VSS VSS nch W=0.8U L=0.24U
M7 TP1 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP1 VDD VDD pch W=2.7U L=0.24U
M10 TP4 TP1 VSS VSS nch W=2.2U L=0.24U
M38 QN Q VSS VSS nch W=2.88U L=0.24U
M30 TP14 Q VDD VDD pch W=1.3U L=0.24U
M33 Q TP13 VDD VDD pch W=6.26U L=0.24U
M23 TP11 TP8 TP12 VSS nch W=2.92U L=0.24U
M13 TP8 CLK DIN VDD pch W=1.3U L=0.24U
M14 DIN TP6 TP8 VSS nch W=0.8U L=0.24U
M25 TP11 CLK TP13 VSS nch W=2.7U L=0.24U
M26 TP13 TP6 TP11 VDD pch W=3U L=0.24U
M15 TP8 CLK TP9 VSS nch W=0.8U L=0.24U
M16 TP9 TP6 TP8 VDD pch W=1.3U L=0.24U
M27 TP14 CLK TP13 VDD pch W=1.3U L=0.24U
M28 TP13 TP6 TP14 VSS nch W=0.8U L=0.24U
M17 TP9 TP2 VDD VDD pch W=1.3U L=0.24U
M21 TP11 TP8 VDD VDD pch W=3.24U L=0.24U
M22 TP11 TP4 VDD VDD pch W=3.24U L=0.24U
M29 TP14 TP4 VDD VDD pch W=1.3U L=0.24U
M37 QN Q VDD VDD pch W=6.2U L=0.24U
M31 TP14 Q TP15 VSS nch W=0.8U L=0.24U
M20 TP10 TP11 VSS VSS nch W=0.8U L=0.24U
M32 TP15 TP4 VSS VSS nch W=0.8U L=0.24U
M24 TP12 TP4 VSS VSS nch W=2.92U L=0.24U
M36 TP16 TP13 VSS VSS nch W=5.26U L=0.24U
M34 Q TP2 VDD VDD pch W=6.26U L=0.24U
M35 Q TP2 TP16 VSS nch W=5.26U L=0.24U
M18 TP9 TP11 VDD VDD pch W=1.3U L=0.24U
M19 TP9 TP2 TP10 VSS nch W=0.8U L=0.24U
M11 TP6 CLK VDD VDD pch W=1.6U L=0.24U
M5 TP2 TP0 TP3 VSS nch W=2.2U L=0.24U
M6 TP3 TP4 VSS VSS nch W=2.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffass1 Q QN SETB CLK DIN
M19 TP7 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 DIN VSS VSS nch W=0.8U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.3U L=0.24U
M23 QN TP8 VDD VDD pch W=3.14U L=0.24U
M11 TP5 TP3 VDD VDD pch W=1.3U L=0.24U
M26 Q QN VSS VSS nch W=1.42U L=0.24U
M5 TP3 CLK TP0 VDD pch W=1.3U L=0.24U
M6 TP0 TP1 TP3 VSS nch W=0.8U L=0.24U
M15 TP5 CLK TP8 VSS nch W=0.96U L=0.24U
M16 TP8 TP1 TP5 VDD pch W=1.4U L=0.24U
M8 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M17 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M18 TP8 TP1 TP7 VSS nch W=0.8U L=0.24U
M25 Q QN VDD VDD pch W=3.02U L=0.24U
M7 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M13 TP5 TP3 TP6 VSS nch W=0.9U L=0.24U
M21 TP7 QN TP9 VSS nch W=0.9U L=0.24U
M24 QN TP8 VSS VSS nch W=1.96U L=0.24U
M12 TP5 SETB VDD VDD pch W=1.3U L=0.24U
M10 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M14 TP6 SETB VSS VSS nch W=0.9U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M20 TP7 QN VDD VDD pch W=1.3U L=0.24U
M22 TP9 SETB VSS VSS nch W=0.9U L=0.24U
M4 TP1 CLK VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffass2 Q QN SETB CLK DIN
M19 TP7 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 DIN VSS VSS nch W=0.8U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.3U L=0.24U
M23 QN TP8 VDD VDD pch W=6.2U L=0.24U
M11 TP5 TP3 VDD VDD pch W=1.84U L=0.24U
M26 Q QN VSS VSS nch W=2.68U L=0.24U
M5 TP3 CLK TP0 VDD pch W=1.3U L=0.24U
M6 TP0 TP1 TP3 VSS nch W=0.8U L=0.24U
M15 TP5 CLK TP8 VSS nch W=1.52U L=0.24U
M16 TP8 TP1 TP5 VDD pch W=1.9U L=0.24U
M8 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M17 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M18 TP8 TP1 TP7 VSS nch W=0.8U L=0.24U
M25 Q QN VDD VDD pch W=6.16U L=0.24U
M7 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M13 TP5 TP3 TP6 VSS nch W=1.48U L=0.24U
M21 TP7 QN TP9 VSS nch W=0.9U L=0.24U
M24 QN TP8 VSS VSS nch W=3.98U L=0.24U
M12 TP5 SETB VDD VDD pch W=1.84U L=0.24U
M10 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M14 TP6 SETB VSS VSS nch W=1.48U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M20 TP7 QN VDD VDD pch W=1.3U L=0.24U
M22 TP9 SETB VSS VSS nch W=0.9U L=0.24U
M4 TP1 CLK VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffcs1 Q QN CLK DIN CLRB
M8 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M9 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M10 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M15 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M17 TP6 CLK TP7 VSS nch W=0.8U L=0.24U
M18 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M23 QN TP7 VDD VDD pch W=3.14U L=0.24U
M24 QN TP7 VSS VSS nch W=2.06U L=0.24U
M11 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M12 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M14 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M19 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M25 Q QN VDD VDD pch W=2.94U L=0.24U
M26 Q QN VSS VSS nch W=1.28U L=0.24U
M16 TP6 TP4 VSS VSS nch W=0.8U L=0.24U
M7 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M22 TP8 QN VSS VSS nch W=0.8U L=0.24U
M20 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M21 TP8 QN VDD VDD pch W=1.3U L=0.24U
M3 TP2 DIN TP1 VSS nch W=0.8U L=0.24U
M13 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M4 TP1 CLRB VSS VSS nch W=0.8U L=0.24U
M2 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M1 TP2 DIN VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffcs2 Q QN CLK DIN CLRB
M8 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M9 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M10 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M15 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M17 TP6 CLK TP7 VSS nch W=1.3U L=0.24U
M18 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M23 QN TP7 VDD VDD pch W=6.24U L=0.24U
M24 QN TP7 VSS VSS nch W=3.98U L=0.24U
M11 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M12 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M14 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M19 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M25 Q QN VDD VDD pch W=5.92U L=0.24U
M26 Q QN VSS VSS nch W=2.66U L=0.24U
M16 TP6 TP4 VSS VSS nch W=1.26U L=0.24U
M7 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M22 TP8 QN VSS VSS nch W=0.8U L=0.24U
M20 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M21 TP8 QN VDD VDD pch W=1.3U L=0.24U
M3 TP2 DIN TP1 VSS nch W=0.8U L=0.24U
M13 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M4 TP1 CLRB VSS VSS nch W=0.8U L=0.24U
M2 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M1 TP2 DIN VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffles1 EB DIN CLK QN Q
M8 N1N80 TP7 VSS VSS nch W=0.8U L=0.24U
M7 N1N80 TP7 VDD VDD pch W=1.3U L=0.24U
M12 TP21 TP1 TP3 VSS nch W=0.8U L=0.24U
M19 TP5 CLK TP6 VSS nch W=0.8U L=0.24U
M20 TP6 TP1 TP5 VDD pch W=1.3U L=0.24U
M26 Q TP6 VSS VSS nch W=2.06U L=0.24U
M13 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M14 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M15 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M16 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M21 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M22 TP6 TP1 TP7 VSS nch W=0.8U L=0.24U
M24 TP7 Q VSS VSS nch W=0.8U L=0.24U
M28 QN Q VSS VSS nch W=1.28U L=0.24U
M18 TP5 TP3 VSS VSS nch W=0.8U L=0.24U
M11 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M17 TP5 TP3 VDD VDD pch W=1.8U L=0.24U
M27 QN Q VDD VDD pch W=2.94U L=0.24U
M25 Q TP6 VDD VDD pch W=3.14U L=0.24U
M9 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M23 TP7 Q VDD VDD pch W=1.3U L=0.24U
M10 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M3 N1N80 EB TP21 VSS nch W=0.8U L=0.24U
M4 TP21 TP20 N1N80 VDD pch W=1.3U L=0.24U
M5 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M6 TP21 EB DIN VDD pch W=1.3U L=0.24U
M1 TP20 EB VDD VDD pch W=1.3U L=0.24U
M2 TP20 EB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffles2 EB DIN CLK QN Q
M8 N1N80 TP7 VSS VSS nch W=0.8U L=0.24U
M7 N1N80 TP7 VDD VDD pch W=1.3U L=0.24U
M12 TP21 TP1 TP3 VSS nch W=0.8U L=0.24U
M19 TP5 CLK TP6 VSS nch W=1.3U L=0.24U
M20 TP6 TP1 TP5 VDD pch W=1.8U L=0.24U
M26 Q TP6 VSS VSS nch W=3.98U L=0.24U
M13 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M14 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M15 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M16 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M21 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M22 TP6 TP1 TP7 VSS nch W=0.8U L=0.24U
M24 TP7 Q VSS VSS nch W=0.8U L=0.24U
M28 QN Q VSS VSS nch W=2.66U L=0.24U
M18 TP5 TP3 VSS VSS nch W=1.26U L=0.24U
M11 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M17 TP5 TP3 VDD VDD pch W=2.78U L=0.24U
M27 QN Q VDD VDD pch W=5.92U L=0.24U
M25 Q TP6 VDD VDD pch W=6.24U L=0.24U
M9 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M23 TP7 Q VDD VDD pch W=1.3U L=0.24U
M10 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M3 N1N80 EB TP21 VSS nch W=0.8U L=0.24U
M4 TP21 TP20 N1N80 VDD pch W=1.3U L=0.24U
M5 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M6 TP21 EB DIN VDD pch W=1.3U L=0.24U
M1 TP20 EB VDD VDD pch W=1.3U L=0.24U
M2 TP20 EB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffs1 QN CLK DIN
M8 DIN TP1 TP3 VSS nch W=0.8U L=0.24U
M15 TP5 CLK TP6 VSS nch W=0.8U L=0.24U
M16 TP6 TP1 TP5 VDD pch W=1.3U L=0.24U
M20 Q TP6 VSS VSS nch W=2.06U L=0.24U
M9 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M10 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M14 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M17 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M18 TP6 TP1 TP7 VSS nch W=0.8U L=0.24U
M21 TP7 Q VDD VDD pch W=1.3U L=0.24U
M22 TP7 Q VSS VSS nch W=0.8U L=0.24U
M24 QN Q VSS VSS nch W=1.28U L=0.24U
M12 TP5 TP3 VSS VSS nch W=0.8U L=0.24U
M7 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M11 TP5 TP3 VDD VDD pch W=1.8U L=0.24U
M23 QN Q VDD VDD pch W=2.94U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M19 Q TP6 VDD VDD pch W=3.14U L=0.24U
M4 TP1 CLK VSS VSS nch W=0.8U L=0.24U
.ENDS

.SUBCKT dffs1 QN Q CLK DIN
M8 DIN TP1 TP3 VSS nch W=0.8U L=0.24U
M15 TP5 CLK TP6 VSS nch W=0.8U L=0.24U
M16 TP6 TP1 TP5 VDD pch W=1.3U L=0.24U
M20 Q TP6 VSS VSS nch W=2.06U L=0.24U
M9 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M10 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M14 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M17 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M18 TP6 TP1 TP7 VSS nch W=0.8U L=0.24U
M21 TP7 Q VDD VDD pch W=1.3U L=0.24U
M22 TP7 Q VSS VSS nch W=0.8U L=0.24U
M24 QN Q VSS VSS nch W=1.28U L=0.24U
M12 TP5 TP3 VSS VSS nch W=0.8U L=0.24U
M7 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M11 TP5 TP3 VDD VDD pch W=1.8U L=0.24U
M23 QN Q VDD VDD pch W=2.94U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M19 Q TP6 VDD VDD pch W=3.14U L=0.24U
M4 TP1 CLK VSS VSS nch W=0.8U L=0.24U
.ENDS

.SUBCKT dffs1 Q CLK DIN
M8 DIN TP1 TP3 VSS nch W=0.8U L=0.24U
M15 TP5 CLK TP6 VSS nch W=0.8U L=0.24U
M16 TP6 TP1 TP5 VDD pch W=1.3U L=0.24U
M20 Q TP6 VSS VSS nch W=2.06U L=0.24U
M9 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M10 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M14 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M17 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M18 TP6 TP1 TP7 VSS nch W=0.8U L=0.24U
M21 TP7 Q VDD VDD pch W=1.3U L=0.24U
M22 TP7 Q VSS VSS nch W=0.8U L=0.24U
M24 QN Q VSS VSS nch W=1.28U L=0.24U
M12 TP5 TP3 VSS VSS nch W=0.8U L=0.24U
M7 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M11 TP5 TP3 VDD VDD pch W=1.8U L=0.24U
M23 QN Q VDD VDD pch W=2.94U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M19 Q TP6 VDD VDD pch W=3.14U L=0.24U
M4 TP1 CLK VSS VSS nch W=0.8U L=0.24U
.ENDS

.SUBCKT dffs2 DIN CLK Q QN
M8 DIN TP1 TP3 VSS nch W=0.8U L=0.24U
M15 TP5 CLK TP6 VSS nch W=1.3U L=0.24U
M16 TP6 TP1 TP5 VDD pch W=1.8U L=0.24U
M20 Q TP6 VSS VSS nch W=3.98U L=0.24U
M9 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M10 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M14 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M17 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M18 TP6 TP1 TP7 VSS nch W=0.8U L=0.24U
M21 TP7 Q VDD VDD pch W=1.3U L=0.24U
M22 TP7 Q VSS VSS nch W=0.8U L=0.24U
M24 QN Q VSS VSS nch W=2.66U L=0.24U
M12 TP5 TP3 VSS VSS nch W=1.26U L=0.24U
M7 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M11 TP5 TP3 VDD VDD pch W=2.76U L=0.24U
M23 QN Q VDD VDD pch W=5.92U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M19 Q TP6 VDD VDD pch W=6.24U L=0.24U
M4 TP1 CLK VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffscs1 DIN SETB CLRB CLK Q OUTB
M11 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M12 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M17 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M19 TP6 CLK TP7 VSS nch W=0.8U L=0.24U
M20 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M25 QN TP7 VDD VDD pch W=3.14U L=0.24U
M26 QN TP7 VSS VSS nch W=2.06U L=0.24U
M13 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M14 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M16 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M21 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M27 Q QN VDD VDD pch W=2.94U L=0.24U
M28 Q QN VSS VSS nch W=1.28U L=0.24U
M18 TP6 TP4 VSS VSS nch W=0.8U L=0.24U
M9 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M10 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M24 TP8 QN VSS VSS nch W=0.8U L=0.24U
M22 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M23 TP8 QN VDD VDD pch W=1.3U L=0.24U
M15 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M4 TP2 DIN TP1 VDD pch W=1.3U L=0.24U
M5 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M6 TP2 CLRB TP9 VSS nch W=0.8U L=0.24U
M7 TP9 DIN VSS VSS nch W=0.8U L=0.24U
M8 TP9 TP0 VSS VSS nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 SETB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffscs2 DIN SETB CLRB CLK Q OUTB
M11 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M12 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M17 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M19 TP6 CLK TP7 VSS nch W=1.3U L=0.24U
M20 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M25 QN TP7 VDD VDD pch W=6.24U L=0.24U
M26 QN TP7 VSS VSS nch W=3.98U L=0.24U
M13 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M14 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M16 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M21 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M27 Q QN VDD VDD pch W=5.92U L=0.24U
M28 Q QN VSS VSS nch W=2.66U L=0.24U
M18 TP6 TP4 VSS VSS nch W=1.26U L=0.24U
M9 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M10 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M24 TP8 QN VSS VSS nch W=0.8U L=0.24U
M22 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M23 TP8 QN VDD VDD pch W=1.3U L=0.24U
M15 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M4 TP2 DIN TP1 VDD pch W=1.3U L=0.24U
M5 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M6 TP2 CLRB TP9 VSS nch W=0.8U L=0.24U
M7 TP9 DIN VSS VSS nch W=0.8U L=0.24U
M8 TP9 TP0 VSS VSS nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 SETB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffss1 SETB DIN CLK QN Q
M5 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M1 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M8 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M9 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M10 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M15 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M17 TP6 CLK TP7 VSS nch W=0.8U L=0.24U
M18 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M23 QN TP7 VDD VDD pch W=3.14U L=0.24U
M24 QN TP7 VSS VSS nch W=2.06U L=0.24U
M11 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M12 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M14 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M19 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M25 Q QN VDD VDD pch W=2.94U L=0.24U
M26 Q QN VSS VSS nch W=1.28U L=0.24U
M16 TP6 TP4 VSS VSS nch W=0.8U L=0.24U
M7 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M22 TP8 QN VSS VSS nch W=0.8U L=0.24U
M2 TP2 DIN TP1 VDD pch W=1.3U L=0.24U
M3 TP2 DIN VSS VSS nch W=0.8U L=0.24U
M4 TP2 TP0 VSS VSS nch W=0.8U L=0.24U
M20 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M21 TP8 QN VDD VDD pch W=1.3U L=0.24U
M13 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M6 TP0 SETB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dffss2 SETB DIN CLK QN Q
M5 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M1 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M8 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M9 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M10 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M15 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M17 TP6 CLK TP7 VSS nch W=1.3U L=0.24U
M18 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M23 QN TP7 VDD VDD pch W=6.24U L=0.24U
M24 QN TP7 VSS VSS nch W=3.98U L=0.24U
M11 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M12 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M14 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M19 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M25 Q QN VDD VDD pch W=5.92U L=0.24U
M26 Q QN VSS VSS nch W=2.66U L=0.24U
M16 TP6 TP4 VSS VSS nch W=1.26U L=0.24U
M7 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M22 TP8 QN VSS VSS nch W=0.8U L=0.24U
M2 TP2 DIN TP1 VDD pch W=1.3U L=0.24U
M3 TP2 DIN VSS VSS nch W=0.8U L=0.24U
M4 TP2 TP0 VSS VSS nch W=0.8U L=0.24U
M20 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M21 TP8 QN VDD VDD pch W=1.3U L=0.24U
M13 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M6 TP0 SETB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s1 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=1.8U L=0.24U
M4 VSS DIN2 Q2 VSS nch W=0.74U L=0.24U
M2 Q1 DIN1 VSS VSS nch W=0.74U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s10 DIN1 DIN2 Q1 Q2
M1 N1N255 DIN1 VDD VDD pch W=9.5U L=0.24U
M2 N1N255 DIN1 VSS VSS nch W=6.8U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=20.28U L=0.24U
M4 N1N266 N1N255 VSS VSS nch W=14.56U L=0.24U
M5 Q1 N1N266 VDD VDD pch W=47.64U L=0.24U
M6 Q1 N1N266 VSS VSS nch W=19.5U L=0.24U
M8 N1N340 DIN2 VSS VSS nch W=6.8U L=0.24U
M7 N1N340 DIN2 VDD VDD pch W=9.5U L=0.24U
M10 N1N347 N1N340 VSS VSS nch W=14.56U L=0.24U
M9 N1N347 N1N340 VDD VDD pch W=20.28U L=0.24U
M12 Q2 N1N347 VSS VSS nch W=19.5U L=0.24U
M11 Q2 N1N347 VDD VDD pch W=47.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s11 DIN1 DIN2 Q1 Q2
M3 N1N255 N1N253 VDD VDD pch W=9U L=0.24U
M4 N1N255 N1N253 VSS VSS nch W=4.5U L=0.24U
M5 N1N266 N1N255 VDD VDD pch W=20U L=0.24U
M6 N1N266 N1N255 VSS VSS nch W=11U L=0.24U
M7 N1N268 N1N266 VDD VDD pch W=40U L=0.24U
M8 N1N268 N1N266 VSS VSS nch W=26U L=0.24U
M1 N1N253 DIN1 VDD VDD pch W=4U L=0.24U
M2 N1N253 DIN1 VSS VSS nch W=2.2U L=0.24U
M9 Q1 N1N268 VDD VDD pch W=84U L=0.24U
M10 Q1 N1N268 VSS VSS nch W=42U L=0.24U
M14 N1N312 N1N299 VSS VSS nch W=4.5U L=0.24U
M13 N1N312 N1N299 VDD VDD pch W=9U L=0.24U
M16 N1N319 N1N312 VSS VSS nch W=11U L=0.24U
M15 N1N319 N1N312 VDD VDD pch W=20U L=0.24U
M18 N1N297 N1N319 VSS VSS nch W=26U L=0.24U
M17 N1N297 N1N319 VDD VDD pch W=40U L=0.24U
M12 N1N299 DIN2 VSS VSS nch W=2.2U L=0.24U
M11 N1N299 DIN2 VDD VDD pch W=4U L=0.24U
M20 Q2 N1N297 VSS VSS nch W=42U L=0.24U
M19 Q2 N1N297 VDD VDD pch W=84U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s12 DIN1 DIN2 Q1 Q2
M3 N1N255 N1N253 VDD VDD pch W=16.5U L=0.24U
M4 N1N255 N1N253 VSS VSS nch W=9.8U L=0.24U
M5 N1N266 N1N255 VDD VDD pch W=36.4U L=0.24U
M6 N1N266 N1N255 VSS VSS nch W=20.6U L=0.24U
M7 N1N268 N1N266 VDD VDD pch W=88.3U L=0.24U
M8 N1N268 N1N266 VSS VSS nch W=50.9U L=0.24U
M1 N1N253 DIN1 VDD VDD pch W=8.3U L=0.24U
M2 N1N253 DIN1 VSS VSS nch W=5U L=0.24U
M9 Q1 N1N268 VDD VDD pch W=180.8U L=0.24U
M10 Q1 N1N268 VSS VSS nch W=78.6U L=0.24U
M14 N1N312 N1N299 VSS VSS nch W=9.8U L=0.24U
M13 N1N312 N1N299 VDD VDD pch W=16.5U L=0.24U
M16 N1N319 N1N312 VSS VSS nch W=20.6U L=0.24U
M15 N1N319 N1N312 VDD VDD pch W=36.4U L=0.24U
M18 N1N297 N1N319 VSS VSS nch W=50.9U L=0.24U
M17 N1N297 N1N319 VDD VDD pch W=88.3U L=0.24U
M12 N1N299 DIN2 VSS VSS nch W=5U L=0.24U
M11 N1N299 DIN2 VDD VDD pch W=8.3U L=0.24U
M20 Q2 N1N297 VSS VSS nch W=78.6U L=0.24U
M19 Q2 N1N297 VDD VDD pch W=180.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s2 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=3.16U L=0.24U
M4 VSS DIN2 Q2 VSS nch W=1.24U L=0.24U
M2 Q1 DIN1 VSS VSS nch W=1.24U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=3.16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s3 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=4.98U L=0.24U
M4 VSS DIN2 Q2 VSS nch W=2.14U L=0.24U
M2 Q1 DIN1 VSS VSS nch W=2.14U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=4.98U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s4 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=5.8U L=0.24U
M4 VSS DIN2 Q2 VSS nch W=2.5U L=0.24U
M2 Q1 DIN1 VSS VSS nch W=2.5U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=5.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s5 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=8.28U L=0.24U
M4 VSS DIN2 Q2 VSS nch W=3.5U L=0.24U
M2 Q1 DIN1 VSS VSS nch W=3.5U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=8.28U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s6 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=10.7U L=0.24U
M4 VSS DIN2 Q2 VSS nch W=4.7U L=0.24U
M2 Q1 DIN1 VSS VSS nch W=4.7U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=10.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s7 DIN1 DIN2 Q1 Q2
M1 N1N255 DIN1 VDD VDD pch W=4.1U L=0.24U
M2 N1N255 DIN1 VSS VSS nch W=1.9U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=5.5U L=0.24U
M4 N1N266 N1N255 VSS VSS nch W=3.1U L=0.24U
M5 Q1 N1N266 VDD VDD pch W=15.2U L=0.24U
M6 Q1 N1N266 VSS VSS nch W=8.5U L=0.24U
M8 N1N340 DIN2 VSS VSS nch W=1.9U L=0.24U
M7 N1N340 DIN2 VDD VDD pch W=4.1U L=0.24U
M10 N1N347 N1N340 VSS VSS nch W=3.1U L=0.24U
M9 N1N347 N1N340 VDD VDD pch W=5.5U L=0.24U
M12 Q2 N1N347 VSS VSS nch W=8.5U L=0.24U
M11 Q2 N1N347 VDD VDD pch W=15.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s8 DIN1 DIN2 Q1 Q2
M1 N1N255 DIN1 VDD VDD pch W=5.6U L=0.24U
M2 N1N255 DIN1 VSS VSS nch W=4U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=12U L=0.24U
M4 N1N266 N1N255 VSS VSS nch W=8.6U L=0.24U
M5 Q1 N1N266 VDD VDD pch W=25.4U L=0.24U
M6 Q1 N1N266 VSS VSS nch W=12.7U L=0.24U
M8 N1N340 DIN2 VSS VSS nch W=4U L=0.24U
M7 N1N340 DIN2 VDD VDD pch W=5.6U L=0.24U
M10 N1N347 N1N340 VSS VSS nch W=8.6U L=0.24U
M9 N1N347 N1N340 VDD VDD pch W=12U L=0.24U
M12 Q2 N1N347 VSS VSS nch W=12.7U L=0.24U
M11 Q2 N1N347 VDD VDD pch W=25.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT di2s9 DIN1 DIN2 Q1 Q2
M1 N1N255 DIN1 VDD VDD pch W=7.3U L=0.24U
M2 N1N255 DIN1 VSS VSS nch W=5.2U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=15.6U L=0.24U
M4 N1N266 N1N255 VSS VSS nch W=11.2U L=0.24U
M5 Q1 N1N266 VDD VDD pch W=35.8U L=0.24U
M6 Q1 N1N266 VSS VSS nch W=15U L=0.24U
M8 N1N340 DIN2 VSS VSS nch W=5.2U L=0.24U
M7 N1N340 DIN2 VDD VDD pch W=7.3U L=0.24U
M10 N1N347 N1N340 VSS VSS nch W=11.2U L=0.24U
M9 N1N347 N1N340 VDD VDD pch W=15.6U L=0.24U
M12 Q2 N1N347 VSS VSS nch W=15U L=0.24U
M11 Q2 N1N347 VDD VDD pch W=35.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dsmxc31s1 Q DIN1 CLK DIN2
M7 N1N280 DIN1 N1N270 VSS nch W=0.6U L=0.24U
M3 N1N261 DIN2 VDD VDD pch W=1.1U L=0.24U
M5 N1N280 N1N276 N1N261 VDD pch W=1.1U L=0.24U
M4 VDD CLK N1N263 VDD pch W=1.1U L=0.24U
M6 N1N263 DIN1 N1N280 VDD pch W=1.1U L=0.24U
M9 N1N270 N1N276 VSS VSS nch W=0.6U L=0.24U
M2 N1N276 CLK VSS VSS nch W=0.6U L=0.24U
M1 N1N276 CLK VDD VDD pch W=1.2U L=0.24U
M8 N1N272 CLK N1N280 VSS nch W=0.6U L=0.24U
M10 VSS DIN2 N1N272 VSS nch W=0.6U L=0.24U
M11 Q N1N280 VDD VDD pch W=1.84U L=0.24U
M12 Q N1N280 VSS VSS nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT dsmxc31s2 Q DIN1 CLK DIN2
M7 N1N280 DIN1 N1N270 VSS nch W=0.8U L=0.24U
M3 N1N261 DIN2 VDD VDD pch W=1.5U L=0.24U
M5 N1N280 N1N276 N1N261 VDD pch W=1.5U L=0.24U
M4 VDD CLK N1N263 VDD pch W=1.5U L=0.24U
M6 N1N263 DIN1 N1N280 VDD pch W=1.5U L=0.24U
M9 N1N270 N1N276 VSS VSS nch W=0.8U L=0.24U
M2 N1N276 CLK VSS VSS nch W=0.6U L=0.24U
M1 N1N276 CLK VDD VDD pch W=1.2U L=0.24U
M8 N1N272 CLK N1N280 VSS nch W=0.8U L=0.24U
M10 VSS DIN2 N1N272 VSS nch W=0.8U L=0.24U
M11 Q N1N280 VDD VDD pch W=2.6U L=0.24U
M12 Q N1N280 VSS VSS nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT fadd1s1 OUTS OUTC AIN BIN CIN
M1 TP9 AIN VDD VDD pch W=1.2U L=0.24U
M2 TP0 BIN TP9 VDD pch W=1.1U L=0.24U
M3 TP0 BIN TP8 VSS nch W=0.8U L=0.24U
M4 TP8 AIN VSS VSS nch W=0.9U L=0.24U
M5 TP10 AIN VDD VDD pch W=1.2U L=0.24U
M6 VDD BIN TP10 VDD pch W=1.2U L=0.24U
M7 TP10 CIN TP0 VDD pch W=1.1U L=0.24U
M8 TP11 CIN TP0 VSS nch W=0.8U L=0.24U
M9 VSS BIN TP11 VSS nch W=0.9U L=0.24U
M10 TP11 AIN VSS VSS nch W=0.9U L=0.24U
M11 TP1 AIN VDD VDD pch W=1.4U L=0.24U
M12 TP3 TP0 TP1 VDD pch W=1.1U L=0.24U
M13 TP3 TP0 TP2 VSS nch W=0.9U L=0.24U
M14 TP2 AIN VSS VSS nch W=0.9U L=0.24U
M15 TP1 BIN VDD VDD pch W=1.4U L=0.24U
M16 VDD CIN TP1 VDD pch W=1.4U L=0.24U
M17 TP2 BIN VSS VSS nch W=0.9U L=0.24U
M18 VSS CIN TP2 VSS nch W=0.9U L=0.24U
M19 VDD AIN TP4 VDD pch W=2.1U L=0.24U
M20 TP4 BIN TP5 VDD pch W=2.1U L=0.24U
M21 TP5 CIN TP3 VDD pch W=2.1U L=0.24U
M22 TP6 CIN TP3 VSS nch W=1.3U L=0.24U
M23 TP7 BIN TP6 VSS nch W=1.3U L=0.24U
M24 VSS AIN TP7 VSS nch W=1.3U L=0.24U
M26 OUTS TP3 VSS VSS nch W=0.9U L=0.24U
M28 OUTC TP0 VSS VSS nch W=1U L=0.24U
M25 OUTS TP3 VDD VDD pch W=1.3U L=0.24U
M27 OUTC TP0 VDD VDD pch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT fadd1s2 OUTS OUTC AIN BIN CIN
M1 TP9 AIN VDD VDD pch W=1.8U L=0.24U
M2 TP0 BIN TP9 VDD pch W=1.7U L=0.24U
M3 TP0 BIN TP8 VSS nch W=1.1U L=0.24U
M4 TP8 AIN VSS VSS nch W=1.2U L=0.24U
M5 TP10 AIN VDD VDD pch W=1.8U L=0.24U
M6 VDD BIN TP10 VDD pch W=1.8U L=0.24U
M7 TP10 CIN TP0 VDD pch W=1.7U L=0.24U
M8 TP11 CIN TP0 VSS nch W=1.1U L=0.24U
M9 VSS BIN TP11 VSS nch W=1.2U L=0.24U
M10 TP11 AIN VSS VSS nch W=1.2U L=0.24U
M11 TP1 AIN VDD VDD pch W=2.1U L=0.24U
M12 TP3 TP0 TP1 VDD pch W=1.66U L=0.24U
M13 TP3 TP0 TP2 VSS nch W=1.16U L=0.24U
M14 TP2 AIN VSS VSS nch W=1.16U L=0.24U
M15 TP1 BIN VDD VDD pch W=2.1U L=0.24U
M16 VDD CIN TP1 VDD pch W=2.1U L=0.24U
M17 TP2 BIN VSS VSS nch W=1.16U L=0.24U
M18 VSS CIN TP2 VSS nch W=1.16U L=0.24U
M19 VDD AIN TP4 VDD pch W=3.16U L=0.24U
M20 TP4 BIN TP5 VDD pch W=3.16U L=0.24U
M21 TP5 CIN TP3 VDD pch W=3.16U L=0.24U
M22 TP6 CIN TP3 VSS nch W=1.74U L=0.24U
M23 TP7 BIN TP6 VSS nch W=1.74U L=0.24U
M24 VSS AIN TP7 VSS nch W=1.74U L=0.24U
M26 OUTS TP3 VSS VSS nch W=1.44U L=0.24U
M28 OUTC TP0 VSS VSS nch W=1.62U L=0.24U
M25 OUTS TP3 VDD VDD pch W=2.1U L=0.24U
M27 OUTC TP0 VDD VDD pch W=2.32U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT fadd1s3 OUTS OUTC AIN BIN CIN
M1 TP9 AIN VDD VDD pch W=2.7U L=0.24U
M2 TP0 BIN TP9 VDD pch W=2.6U L=0.24U
M3 TP0 BIN TP8 VSS nch W=1.6U L=0.24U
M4 TP8 AIN VSS VSS nch W=1.7U L=0.24U
M5 TP10 AIN VDD VDD pch W=2.7U L=0.24U
M6 VDD BIN TP10 VDD pch W=2.7U L=0.24U
M7 TP10 CIN TP0 VDD pch W=2.6U L=0.24U
M8 TP11 CIN TP0 VSS nch W=1.6U L=0.24U
M9 VSS BIN TP11 VSS nch W=1.7U L=0.24U
M10 TP11 AIN VSS VSS nch W=1.7U L=0.24U
M11 TP1 AIN VDD VDD pch W=2.9U L=0.24U
M12 TP3 TP0 TP1 VDD pch W=2.8U L=0.24U
M13 TP3 TP0 TP2 VSS nch W=1.52U L=0.24U
M14 TP2 AIN VSS VSS nch W=1.52U L=0.24U
M15 TP1 BIN VDD VDD pch W=2.9U L=0.24U
M16 VDD CIN TP1 VDD pch W=2.9U L=0.24U
M17 TP2 BIN VSS VSS nch W=1.52U L=0.24U
M18 VSS CIN TP2 VSS nch W=1.52U L=0.24U
M19 VDD AIN TP4 VDD pch W=4.4U L=0.24U
M20 TP4 BIN TP5 VDD pch W=4.4U L=0.24U
M21 TP5 CIN TP3 VDD pch W=4.3U L=0.24U
M22 TP6 CIN TP3 VSS nch W=2.26U L=0.24U
M23 TP7 BIN TP6 VSS nch W=2.26U L=0.24U
M24 VSS AIN TP7 VSS nch W=2.26U L=0.24U
M26 OUTS TP3 VSS VSS nch W=3.1U L=0.24U
M28 OUTC TP0 VSS VSS nch W=3.4U L=0.24U
M25 OUTS TP3 VDD VDD pch W=4.2U L=0.24U
M27 OUTC TP0 VDD VDD pch W=4.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT faddpgs1 AIN BIN CIN OUTG OUTP OUTS
M24 OUTG N1N525 VSS VSS nch W=0.9U L=0.24U
M23 OUTG N1N525 VDD VDD pch W=1.9U L=0.24U
M19 N1N525 AIN N1N553 VSS nch W=0.8U L=0.24U
M17 VDD AIN N1N525 VDD pch W=0.9U L=0.24U
M18 N1N525 BIN VDD VDD pch W=0.9U L=0.24U
M20 N1N553 BIN VSS VSS nch W=0.8U L=0.24U
M5 N1N515 AIN BIN VDD pch W=1.2U L=0.24U
M6 BIN N1N569 N1N515 VSS nch W=0.8U L=0.24U
M1 N1N569 AIN VDD VDD pch W=1.5U L=0.24U
M8 BIN AIN N1N623 VSS nch W=0.8U L=0.24U
M3 N1N572 CIN VDD VDD pch W=1.5U L=0.24U
M4 N1N572 CIN VSS VSS nch W=0.7U L=0.24U
M2 N1N569 AIN VSS VSS nch W=0.7U L=0.24U
M7 N1N623 N1N569 BIN VDD pch W=1.2U L=0.24U
M13 N1N515 BIN AIN VDD pch W=1.6U L=0.24U
M14 N1N515 BIN N1N569 VSS nch W=0.7U L=0.24U
M16 N1N623 BIN AIN VSS nch W=0.7U L=0.24U
M15 N1N623 BIN N1N569 VDD pch W=1.6U L=0.24U
M9 N1N693 N1N515 N1N572 VDD pch W=1.2U L=0.24U
M10 N1N572 N1N623 N1N693 VSS nch W=0.7U L=0.24U
M11 N1N693 N1N623 CIN VDD pch W=1.2U L=0.24U
M12 CIN N1N515 N1N693 VSS nch W=0.7U L=0.24U
M21 OUTS N1N693 VDD VDD pch W=1.4U L=0.24U
M22 OUTS N1N693 VSS VSS nch W=0.9U L=0.24U
M25 OUTP N1N623 VDD VDD pch W=1.9U L=0.24U
M26 OUTP N1N623 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT faddpgs2 AIN BIN CIN OUTG OUTP OUTS
M24 OUTG N1N525 VSS VSS nch W=1.1U L=0.24U
M23 OUTG N1N525 VDD VDD pch W=2.47U L=0.24U
M19 N1N525 AIN N1N553 VSS nch W=0.96U L=0.24U
M17 VDD AIN N1N525 VDD pch W=1.16U L=0.24U
M18 N1N525 BIN VDD VDD pch W=1.16U L=0.24U
M20 N1N553 BIN VSS VSS nch W=0.96U L=0.24U
M5 N1N515 AIN BIN VDD pch W=1.56U L=0.24U
M6 BIN N1N569 N1N515 VSS nch W=1U L=0.24U
M1 N1N569 AIN VDD VDD pch W=1.96U L=0.24U
M8 BIN AIN N1N623 VSS nch W=1U L=0.24U
M3 N1N572 CIN VDD VDD pch W=1.96U L=0.24U
M4 N1N572 CIN VSS VSS nch W=0.92U L=0.24U
M2 N1N569 AIN VSS VSS nch W=0.92U L=0.24U
M7 N1N623 N1N569 BIN VDD pch W=1.5U L=0.24U
M13 N1N515 BIN AIN VDD pch W=1.92U L=0.24U
M14 N1N515 BIN N1N569 VSS nch W=0.84U L=0.24U
M16 N1N623 BIN AIN VSS nch W=0.84U L=0.24U
M15 N1N623 BIN N1N569 VDD pch W=1.92U L=0.24U
M9 N1N693 N1N515 N1N572 VDD pch W=1.56U L=0.24U
M10 N1N572 N1N623 N1N693 VSS nch W=0.84U L=0.24U
M11 N1N693 N1N623 CIN VDD pch W=1.56U L=0.24U
M12 CIN N1N515 N1N693 VSS nch W=0.84U L=0.24U
M21 OUTS N1N693 VDD VDD pch W=1.82U L=0.24U
M22 OUTS N1N693 VSS VSS nch W=1.26U L=0.24U
M25 OUTP N1N623 VDD VDD pch W=2.47U L=0.24U
M26 OUTP N1N623 VSS VSS nch W=1.68U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT faddpgs3 AIN BIN CIN OUTG OUTP OUTS
M24 OUTG N1N525 VSS VSS nch W=1.85U L=0.24U
M23 OUTG N1N525 VDD VDD pch W=3.72U L=0.24U
M19 N1N525 AIN N1N553 VSS nch W=1.44U L=0.24U
M17 VDD AIN N1N525 VDD pch W=1.74U L=0.24U
M18 N1N525 BIN VDD VDD pch W=1.74U L=0.24U
M20 N1N553 BIN VSS VSS nch W=1.44U L=0.24U
M5 N1N515 AIN BIN VDD pch W=2.2U L=0.24U
M6 BIN N1N569 N1N515 VSS nch W=1.6U L=0.24U
M1 N1N569 AIN VDD VDD pch W=2.94U L=0.24U
M8 BIN AIN N1N623 VSS nch W=1.6U L=0.24U
M3 N1N572 CIN VDD VDD pch W=2.34U L=0.24U
M4 N1N572 CIN VSS VSS nch W=1.18U L=0.24U
M2 N1N569 AIN VSS VSS nch W=1.38U L=0.24U
M7 N1N623 N1N569 BIN VDD pch W=2.2U L=0.24U
M13 N1N515 BIN AIN VDD pch W=2.92U L=0.24U
M14 N1N515 BIN N1N569 VSS nch W=1.3U L=0.24U
M16 N1N623 BIN AIN VSS nch W=1.3U L=0.24U
M15 N1N623 BIN N1N569 VDD pch W=2.92U L=0.24U
M9 N1N693 N1N515 N1N572 VDD pch W=2.34U L=0.24U
M10 N1N572 N1N623 N1N693 VSS nch W=1.26U L=0.24U
M11 N1N693 N1N623 CIN VDD pch W=2.34U L=0.24U
M12 CIN N1N515 N1N693 VSS nch W=1.26U L=0.24U
M21 OUTS N1N693 VDD VDD pch W=2.7U L=0.24U
M22 OUTS N1N693 VSS VSS nch W=2.1U L=0.24U
M25 OUTP N1N623 VDD VDD pch W=3.71U L=0.24U
M26 OUTP N1N623 VSS VSS nch W=2.72U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT hadd1s1 AIN BIN OUTS OUTC
M10 VSS BIN N1N458 VSS nch W=0.7U L=0.24U
M7 N1N450 BIN N1N452 VDD pch W=1.6U L=0.24U
M1 N1N439 AIN VDD VDD pch W=0.8U L=0.24U
M5 N1N452 N1N439 VDD VDD pch W=0.8U L=0.24U
M2 VDD BIN N1N439 VDD pch W=0.8U L=0.24U
M6 VDD AIN N1N450 VDD pch W=1.6U L=0.24U
M3 N1N439 AIN N1N443 VSS nch W=0.76U L=0.24U
M4 N1N443 BIN VSS VSS nch W=0.76U L=0.24U
M8 N1N452 N1N439 N1N458 VSS nch W=0.7U L=0.24U
M9 N1N458 AIN VSS VSS nch W=0.7U L=0.24U
M12 OUTS N1N452 VSS VSS nch W=1.16U L=0.24U
M14 OUTC N1N439 VSS VSS nch W=1.4U L=0.24U
M13 OUTC N1N439 VDD VDD pch W=2U L=0.24U
M11 OUTS N1N452 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT hadd1s2 AIN BIN OUTS OUTC
M10 VSS BIN N1N458 VSS nch W=1.1U L=0.24U
M7 N1N450 BIN N1N452 VDD pch W=2.68U L=0.24U
M1 N1N439 AIN VDD VDD pch W=1.4U L=0.24U
M5 N1N452 N1N439 VDD VDD pch W=1.34U L=0.24U
M2 VDD BIN N1N439 VDD pch W=1.4U L=0.24U
M6 VDD AIN N1N450 VDD pch W=2.68U L=0.24U
M3 N1N439 AIN N1N443 VSS nch W=1.14U L=0.24U
M4 N1N443 BIN VSS VSS nch W=1.14U L=0.24U
M8 N1N452 N1N439 N1N458 VSS nch W=1.1U L=0.24U
M9 N1N458 AIN VSS VSS nch W=1.1U L=0.24U
M12 OUTS N1N452 VSS VSS nch W=1.74U L=0.24U
M14 OUTC N1N439 VSS VSS nch W=2.1U L=0.24U
M13 OUTC N1N439 VDD VDD pch W=3U L=0.24U
M11 OUTS N1N452 VDD VDD pch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT hadd1s3 AIN BIN OUTS OUTC
M10 VSS BIN N1N458 VSS nch W=2.2U L=0.24U
M7 N1N450 BIN N1N452 VDD pch W=5.6U L=0.24U
M1 N1N439 AIN VDD VDD pch W=2.9U L=0.24U
M5 N1N452 N1N439 VDD VDD pch W=2.8U L=0.24U
M2 VDD BIN N1N439 VDD pch W=2.9U L=0.24U
M6 VDD AIN N1N450 VDD pch W=5.6U L=0.24U
M3 N1N439 AIN N1N443 VSS nch W=2.28U L=0.24U
M4 N1N443 BIN VSS VSS nch W=2.28U L=0.24U
M8 N1N452 N1N439 N1N458 VSS nch W=2.2U L=0.24U
M9 N1N458 AIN VSS VSS nch W=2.2U L=0.24U
M12 OUTS N1N452 VSS VSS nch W=3.48U L=0.24U
M14 OUTC N1N439 VSS VSS nch W=4.4U L=0.24U
M13 OUTC N1N439 VDD VDD pch W=6U L=0.24U
M11 OUTS N1N452 VDD VDD pch W=5.94U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT hi1s1 Q DIN
M2 Q DIN VSS VSS nch W=0.6U L=0.8U
M1 Q DIN VDD VDD pch W=1U L=0.3U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT hib1s1 Q DIN
M2 Q VSS TP0 VDD pch W=4U L=0.24U
M3 Q VDD TP1 VSS nch W=2U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.9U L=0.4U
M4 TP1 DIN VSS VSS nch W=0.76U L=0.7U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT hnb1s1 Q DIN
M5 Q VDD TP2 VSS nch W=2U L=0.24U
M4 Q VSS TP1 VDD pch W=4U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.6U L=0.24U
M2 TP0 DIN VSS VSS nch W=0.7U L=0.24U
M3 TP1 TP0 VDD VDD pch W=1.9U L=0.4U
M6 TP2 TP0 VSS VSS nch W=0.76U L=0.7U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s1 Q DIN
M1 Q DIN VDD VDD pch W=2U L=0.24U
M2 Q DIN VSS VSS nch W=0.82U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s10 DIN Q
M1 N1N255 DIN VDD VDD pch W=10.5U L=0.24U
M2 N1N255 DIN VSS VSS nch W=6.8U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=21.8U L=0.24U
M4 N1N266 N1N255 VSS VSS nch W=13.6U L=0.24U
M5 Q N1N266 VDD VDD pch W=51.6U L=0.24U
M6 Q N1N266 VSS VSS nch W=20.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s11 DIN Q
M3 N1N255 N1N253 VDD VDD pch W=9U L=0.24U
M4 N1N255 N1N253 VSS VSS nch W=4.5U L=0.24U
M5 N1N266 N1N255 VDD VDD pch W=20U L=0.24U
M6 N1N266 N1N255 VSS VSS nch W=11U L=0.24U
M7 N1N268 N1N266 VDD VDD pch W=40U L=0.24U
M8 N1N268 N1N266 VSS VSS nch W=26U L=0.24U
M1 N1N253 DIN VDD VDD pch W=4U L=0.24U
M2 N1N253 DIN VSS VSS nch W=2.2U L=0.24U
M9 Q N1N268 VDD VDD pch W=84U L=0.24U
M10 Q N1N268 VSS VSS nch W=42U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s12 DIN Q
M3 N1N255 N1N253 VDD VDD pch W=16.5U L=0.24U
M4 N1N255 N1N253 VSS VSS nch W=9.8U L=0.24U
M5 N1N266 N1N255 VDD VDD pch W=36.4U L=0.24U
M6 N1N266 N1N255 VSS VSS nch W=20.6U L=0.24U
M7 N1N268 N1N266 VDD VDD pch W=88.3U L=0.24U
M8 N1N268 N1N266 VSS VSS nch W=50.9U L=0.24U
M1 N1N253 DIN VDD VDD pch W=8.3U L=0.24U
M2 N1N253 DIN VSS VSS nch W=5U L=0.24U
M9 Q N1N268 VDD VDD pch W=180.8U L=0.24U
M10 Q N1N268 VSS VSS nch W=78.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s2 Q DIN
M1 Q DIN VDD VDD pch W=3.5U L=0.24U
M2 Q DIN VSS VSS nch W=1.38U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s3 Q DIN
M1 Q DIN VDD VDD pch W=6.22U L=0.24U
M2 Q DIN VSS VSS nch W=2.68U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s4 Q DIN
M1 Q DIN VDD VDD pch W=7.8U L=0.24U
M2 Q DIN VSS VSS nch W=3.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s5 Q DIN
M1 Q DIN VDD VDD pch W=9.54U L=0.24U
M2 Q DIN VSS VSS nch W=4.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s6 Q DIN
M1 Q DIN VDD VDD pch W=12.6U L=0.24U
M2 Q DIN VSS VSS nch W=5.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s7 Q DIN
M1 N1N255 DIN VDD VDD pch W=4.5U L=0.24U
M2 N1N255 DIN VSS VSS nch W=2.1U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=5.3U L=0.24U
M4 N1N266 N1N255 VSS VSS nch W=4U L=0.24U
M5 Q N1N266 VDD VDD pch W=16.5U L=0.24U
M6 Q N1N266 VSS VSS nch W=9.52U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s8 DIN Q
M1 N1N255 DIN VDD VDD pch W=6.2U L=0.24U
M2 N1N255 DIN VSS VSS nch W=4.5U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=13.5U L=0.24U
M4 N1N266 N1N255 VSS VSS nch W=9.5U L=0.24U
M5 Q N1N266 VDD VDD pch W=28.5U L=0.24U
M6 Q N1N266 VSS VSS nch W=14.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT i1s9 Q DIN
M1 N1N255 DIN VDD VDD pch W=7.3U L=0.24U
M2 N1N255 DIN VSS VSS nch W=5.2U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=15.6U L=0.24U
M4 N1N266 N1N255 VSS VSS nch W=11.2U L=0.24U
M5 Q N1N266 VDD VDD pch W=35.8U L=0.24U
M6 Q N1N266 VSS VSS nch W=15U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s1 Q DIN
M2 Q DIN VSS VSS nch W=1.2U L=0.24U
M1 Q DIN VDD VDD pch W=2.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s10 DIN Q
M2 Q DIN VSS VSS nch W=11.1U L=0.24U
M1 Q DIN VDD VDD pch W=25U L=0.24U
M13 Q DIN VDD VDD pch W=25U L=0.24U
M14 Q DIN VSS VSS nch W=11.1U L=0.24U
M3 Q DIN VDD VDD pch W=25U L=0.24U
M5 Q DIN VDD VDD pch W=25U L=0.24U
M7 Q DIN VDD VDD pch W=25U L=0.24U
M9 Q DIN VDD VDD pch W=25U L=0.24U
M11 Q DIN VDD VDD pch W=25U L=0.24U
M4 Q DIN VSS VSS nch W=11.1U L=0.24U
M6 Q DIN VSS VSS nch W=11.1U L=0.24U
M8 Q DIN VSS VSS nch W=11.1U L=0.24U
M10 Q DIN VSS VSS nch W=11.1U L=0.24U
M12 Q DIN VSS VSS nch W=11.1U L=0.24U
M15 Q DIN VDD VDD pch W=25U L=0.24U
M17 Q DIN VDD VDD pch W=25U L=0.24U
M19 Q DIN VDD VDD pch W=25U L=0.24U
M16 Q DIN VSS VSS nch W=11.1U L=0.24U
M18 Q DIN VSS VSS nch W=11.1U L=0.24U
M20 Q DIN VSS VSS nch W=11.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s11 DIN Q
M2 Q DIN VSS VSS nch W=23U L=0.24U
M1 Q DIN VDD VDD pch W=50U L=0.24U
M13 Q DIN VDD VDD pch W=50U L=0.24U
M14 Q DIN VSS VSS nch W=23U L=0.24U
M3 Q DIN VDD VDD pch W=50U L=0.24U
M5 Q DIN VDD VDD pch W=50U L=0.24U
M7 Q DIN VDD VDD pch W=50U L=0.24U
M9 Q DIN VDD VDD pch W=50U L=0.24U
M11 Q DIN VDD VDD pch W=50U L=0.24U
M4 Q DIN VSS VSS nch W=23U L=0.24U
M6 Q DIN VSS VSS nch W=23U L=0.24U
M8 Q DIN VSS VSS nch W=23U L=0.24U
M10 Q DIN VSS VSS nch W=23U L=0.24U
M12 Q DIN VSS VSS nch W=23U L=0.24U
M15 Q DIN VDD VDD pch W=50U L=0.24U
M17 Q DIN VDD VDD pch W=50U L=0.24U
M19 Q DIN VDD VDD pch W=50U L=0.24U
M16 Q DIN VSS VSS nch W=23U L=0.24U
M18 Q DIN VSS VSS nch W=23U L=0.24U
M20 Q DIN VSS VSS nch W=23U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s12 DIN Q
M2 Q DIN VSS VSS nch W=47U L=0.24U
M1 Q DIN VDD VDD pch W=101U L=0.24U
M13 Q DIN VDD VDD pch W=101U L=0.24U
M14 Q DIN VSS VSS nch W=47U L=0.24U
M3 Q DIN VDD VDD pch W=101U L=0.24U
M5 Q DIN VDD VDD pch W=101U L=0.24U
M7 Q DIN VDD VDD pch W=101U L=0.24U
M9 Q DIN VDD VDD pch W=101U L=0.24U
M11 Q DIN VDD VDD pch W=101U L=0.24U
M4 Q DIN VSS VSS nch W=47U L=0.24U
M6 Q DIN VSS VSS nch W=47U L=0.24U
M8 Q DIN VSS VSS nch W=47U L=0.24U
M10 Q DIN VSS VSS nch W=47U L=0.24U
M12 Q DIN VSS VSS nch W=47U L=0.24U
M15 Q DIN VDD VDD pch W=101U L=0.24U
M17 Q DIN VDD VDD pch W=101U L=0.24U
M19 Q DIN VDD VDD pch W=101U L=0.24U
M16 Q DIN VSS VSS nch W=47U L=0.24U
M18 Q DIN VSS VSS nch W=47U L=0.24U
M20 Q DIN VSS VSS nch W=47U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s2 Q DIN
M2 Q DIN VSS VSS nch W=1.2U L=0.24U
M1 Q DIN VDD VDD pch W=2.9U L=0.24U
M4 Q DIN VSS VSS nch W=1.2U L=0.24U
M3 Q DIN VDD VDD pch W=2.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s3 Q DIN
M2 Q DIN VSS VSS nch W=1.2U L=0.24U
M1 Q DIN VDD VDD pch W=2.9U L=0.24U
M4 Q DIN VSS VSS nch W=1.2U L=0.24U
M3 Q DIN VDD VDD pch W=2.9U L=0.24U
M6 Q DIN VSS VSS nch W=1.2U L=0.24U
M5 Q DIN VDD VDD pch W=2.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s4 Q DIN
M2 Q DIN VSS VSS nch W=1.1U L=0.24U
M1 Q DIN VDD VDD pch W=2.6U L=0.24U
M4 Q DIN VSS VSS nch W=1.1U L=0.24U
M3 Q DIN VDD VDD pch W=2.6U L=0.24U
M6 Q DIN VSS VSS nch W=1.1U L=0.24U
M5 Q DIN VDD VDD pch W=2.6U L=0.24U
M7 Q DIN VDD VDD pch W=2.6U L=0.24U
M8 Q DIN VSS VSS nch W=1.1U L=0.24U
M10 Q DIN VSS VSS nch W=1.1U L=0.24U
M9 Q DIN VDD VDD pch W=2.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s5 Q DIN
M2 Q DIN VSS VSS nch W=1.1U L=0.24U
M1 Q DIN VDD VDD pch W=2.5U L=0.24U
M4 Q DIN VSS VSS nch W=1.1U L=0.24U
M3 Q DIN VDD VDD pch W=2.5U L=0.24U
M6 Q DIN VSS VSS nch W=1.1U L=0.24U
M5 Q DIN VDD VDD pch W=2.5U L=0.24U
M7 Q DIN VDD VDD pch W=2.5U L=0.24U
M8 Q DIN VSS VSS nch W=1.1U L=0.24U
M10 Q DIN VSS VSS nch W=1.1U L=0.24U
M9 Q DIN VDD VDD pch W=2.5U L=0.24U
M12 Q DIN VSS VSS nch W=1.1U L=0.24U
M11 Q DIN VDD VDD pch W=2.5U L=0.24U
M14 Q DIN VSS VSS nch W=1.1U L=0.24U
M13 Q DIN VDD VDD pch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s6 DIN Q
M2 Q DIN VSS VSS nch W=1.1U L=0.24U
M1 Q DIN VDD VDD pch W=2.5U L=0.24U
M4 Q DIN VSS VSS nch W=1.1U L=0.24U
M3 Q DIN VDD VDD pch W=2.5U L=0.24U
M6 Q DIN VSS VSS nch W=1.1U L=0.24U
M5 Q DIN VDD VDD pch W=2.5U L=0.24U
M7 Q DIN VDD VDD pch W=2.5U L=0.24U
M8 Q DIN VSS VSS nch W=1.1U L=0.24U
M10 Q DIN VSS VSS nch W=1.1U L=0.24U
M9 Q DIN VDD VDD pch W=2.5U L=0.24U
M12 Q DIN VSS VSS nch W=1.1U L=0.24U
M11 Q DIN VDD VDD pch W=2.5U L=0.24U
M19 Q DIN VDD VDD pch W=2.5U L=0.24U
M13 Q DIN VDD VDD pch W=2.5U L=0.24U
M16 Q DIN VSS VSS nch W=1.1U L=0.24U
M18 Q DIN VSS VSS nch W=1.1U L=0.24U
M17 Q DIN VDD VDD pch W=2.5U L=0.24U
M14 Q DIN VSS VSS nch W=1.1U L=0.24U
M15 Q DIN VDD VDD pch W=2.5U L=0.24U
M20 Q DIN VSS VSS nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s7 DIN Q
M2 Q DIN VSS VSS nch W=1.8U L=0.24U
M1 Q DIN VDD VDD pch W=4.2U L=0.24U
M13 Q DIN VDD VDD pch W=4.2U L=0.24U
M14 Q DIN VSS VSS nch W=1.8U L=0.24U
M3 Q DIN VDD VDD pch W=4.2U L=0.24U
M5 Q DIN VDD VDD pch W=4.2U L=0.24U
M7 Q DIN VDD VDD pch W=4.2U L=0.24U
M9 Q DIN VDD VDD pch W=4.2U L=0.24U
M11 Q DIN VDD VDD pch W=4.2U L=0.24U
M4 Q DIN VSS VSS nch W=1.8U L=0.24U
M6 Q DIN VSS VSS nch W=1.8U L=0.24U
M8 Q DIN VSS VSS nch W=1.8U L=0.24U
M10 Q DIN VSS VSS nch W=1.8U L=0.24U
M12 Q DIN VSS VSS nch W=1.8U L=0.24U
M15 Q DIN VDD VDD pch W=4.2U L=0.24U
M17 Q DIN VDD VDD pch W=4.2U L=0.24U
M19 Q DIN VDD VDD pch W=4.2U L=0.24U
M16 Q DIN VSS VSS nch W=1.8U L=0.24U
M18 Q DIN VSS VSS nch W=1.8U L=0.24U
M20 Q DIN VSS VSS nch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s8 DIN Q
M2 Q DIN VSS VSS nch W=3.2U L=0.24U
M1 Q DIN VDD VDD pch W=7.5U L=0.24U
M13 Q DIN VDD VDD pch W=7.5U L=0.24U
M14 Q DIN VSS VSS nch W=3.2U L=0.24U
M3 Q DIN VDD VDD pch W=7.5U L=0.24U
M5 Q DIN VDD VDD pch W=7.5U L=0.24U
M7 Q DIN VDD VDD pch W=7.5U L=0.24U
M9 Q DIN VDD VDD pch W=7.5U L=0.24U
M11 Q DIN VDD VDD pch W=7.5U L=0.24U
M4 Q DIN VSS VSS nch W=3.2U L=0.24U
M6 Q DIN VSS VSS nch W=3.2U L=0.24U
M8 Q DIN VSS VSS nch W=3.2U L=0.24U
M10 Q DIN VSS VSS nch W=3.2U L=0.24U
M12 Q DIN VSS VSS nch W=3.2U L=0.24U
M15 Q DIN VDD VDD pch W=7.5U L=0.24U
M17 Q DIN VDD VDD pch W=7.5U L=0.24U
M19 Q DIN VDD VDD pch W=7.5U L=0.24U
M16 Q DIN VSS VSS nch W=3.2U L=0.24U
M18 Q DIN VSS VSS nch W=3.2U L=0.24U
M20 Q DIN VSS VSS nch W=3.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ib1s9 DIN Q
M2 Q DIN VSS VSS nch W=6U L=0.24U
M1 Q DIN VDD VDD pch W=14U L=0.24U
M13 Q DIN VDD VDD pch W=14U L=0.24U
M14 Q DIN VSS VSS nch W=6U L=0.24U
M3 Q DIN VDD VDD pch W=14U L=0.24U
M5 Q DIN VDD VDD pch W=14U L=0.24U
M7 Q DIN VDD VDD pch W=14U L=0.24U
M9 Q DIN VDD VDD pch W=14U L=0.24U
M11 Q DIN VDD VDD pch W=14U L=0.24U
M4 Q DIN VSS VSS nch W=6U L=0.24U
M6 Q DIN VSS VSS nch W=6U L=0.24U
M8 Q DIN VSS VSS nch W=6U L=0.24U
M10 Q DIN VSS VSS nch W=6U L=0.24U
M12 Q DIN VSS VSS nch W=6U L=0.24U
M15 Q DIN VDD VDD pch W=14U L=0.24U
M17 Q DIN VDD VDD pch W=14U L=0.24U
M19 Q DIN VDD VDD pch W=14U L=0.24U
M16 Q DIN VSS VSS nch W=6U L=0.24U
M18 Q DIN VSS VSS nch W=6U L=0.24U
M20 Q DIN VSS VSS nch W=6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lclks1 DIN CLK QN Q
M10 QN TP1 VSS VSS nch W=1.56U L=0.24U
M4 TP1 TP0 DIN VDD pch W=1.8U L=0.24U
M3 DIN CLK TP1 VSS nch W=0.8U L=0.24U
M8 TP2 QN VSS VSS nch W=0.8U L=0.24U
M11 Q QN VDD VDD pch W=2.92U L=0.24U
M12 Q QN VSS VSS nch W=1.34U L=0.24U
M9 QN TP1 VDD VDD pch W=2.92U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M6 TP1 TP0 TP2 VSS nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT holdLatch Q DIN1 DIN2
M10 QN TP1 VSS VSS nch W=1.56U L=0.24U
M4 TP1 TP0 DIN2 VDD pch W=1.8U L=0.24U
M3 DIN2 CLK TP1 VSS nch W=0.8U L=0.24U
M8 TP2 QN VSS VSS nch W=0.8U L=0.24U
M11 Q QN VDD VDD pch W=2.92U L=0.24U
M12 Q QN VSS VSS nch W=1.34U L=0.24U
M9 QN TP1 VDD VDD pch W=2.92U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M6 TP1 TP0 TP2 VSS nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lclks2 DIN CLK QN Q
M10 QN TP1 VSS VSS nch W=3.38U L=0.24U
M4 TP1 TP0 DIN VDD pch W=2.2U L=0.24U
M3 DIN CLK TP1 VSS nch W=1U L=0.24U
M8 TP2 QN VSS VSS nch W=0.8U L=0.24U
M11 Q QN VDD VDD pch W=6.06U L=0.24U
M12 Q QN VSS VSS nch W=2.88U L=0.24U
M9 QN TP1 VDD VDD pch W=6.16U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M6 TP1 TP0 TP2 VSS nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lcs1 CLRB DIN CLK QN Q
M9 QN TP1 VDD VDD pch W=3.1U L=0.24U
M10 QN CLRB VDD VDD pch W=3.1U L=0.24U
M12 TP3 CLRB VSS VSS nch W=2.56U L=0.24U
M11 QN TP1 TP3 VSS nch W=2.56U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK VSS VSS nch W=0.8U L=0.24U
M4 TP1 TP0 DIN VDD pch W=1.88U L=0.24U
M3 DIN CLK TP1 VSS nch W=0.84U L=0.24U
M6 TP1 TP0 TP2 VSS nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M8 TP2 QN VSS VSS nch W=0.8U L=0.24U
M13 Q QN VDD VDD pch W=3.16U L=0.24U
M14 Q QN VSS VSS nch W=1.48U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lcs2 CLRB DIN CLK QN Q
M9 QN TP1 VDD VDD pch W=5.6U L=0.24U
M10 QN CLRB VDD VDD pch W=5.6U L=0.24U
M12 TP3 CLRB VSS VSS nch W=5.1U L=0.24U
M11 QN TP1 TP3 VSS nch W=5.1U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK VSS VSS nch W=0.8U L=0.24U
M4 TP1 TP0 DIN VDD pch W=2.38U L=0.24U
M3 DIN CLK TP1 VSS nch W=1.56U L=0.24U
M6 TP1 TP0 TP2 VSS nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M8 TP2 QN VSS VSS nch W=0.8U L=0.24U
M13 Q QN VDD VDD pch W=6.36U L=0.24U
M14 Q QN VSS VSS nch W=2.94U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lnnds1 Q QN SIN RIN
M1 Q SIN  VDD  VDD P  W=1.56u   L=0.24U
M2 Q QN VDD  VDD P  W=1.56u   L=0.24U
M3 Q QN TP0  VSS   N  W=1.02U   L=0.24U
M4 TP0 SIN  VSS    VSS   N  W=1.02u   L=0.24U
M5 VDD Q  QN VDD P  W=1.56u   L=0.24U
M6 VDD RIN  QN VDD P  W=1.56u   L=0.24U
M7 TP1 Q  QN VSS   N  W=1.02U   L=0.24U
M8 VSS   RIN  TP1  VSS   N  W=1.02u   L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lnnds2 Q QN SIN RIN
M1 Q SIN  VDD  VDD P  W=3.16u  L=0.24U
M2 Q QN VDD  VDD P  W=3.16u  L=0.24U
M3 Q QN TP0  VSS   N  W=2.06U  L=0.24U
M4 TP0 SIN  VSS    VSS   N  W=2.06u  L=0.24U
M5 VDD Q  QN VDD P  W=3.16u  L=0.24U
M6 VDD RIN  QN VDD P  W=3.16u  L=0.24U
M7 TP1 Q  QN VSS   N  W=2.06U  L=0.24U
M8 VSS   RIN  TP1  VSS   N  W=2.06u  L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lnors1 Q QN RIN SIN
M1  TP0   SIN   VDD    VDD  pch W=3.54u    L=0.24U
M2  QN  Q   TP0    VDD  pch W=3.54u    L=0.24U
M3  QN  SIN   VSS      VSS    nch W=0.9u     L=0.24U
M4  VSS     Q   QN   VSS    nch W=0.9u     L=0.24U
M5  VDD  RIN    TP1    VDD  pch W=3.54u    L=0.24U
M6  TP1  QN   Q    VDD  pch W=3.54u    L=0.24U
M7  Q  QN   VSS      VSS    nch W=0.9u     L=0.24U
M8  VSS    RIN    Q    VSS    nch W=0.9u     L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lnors2 Q QN RIN SIN
M1  TP0   SIN   VDD    VDD  pch W=7.18u    L=0.24U
M2  QN  Q   TP0    VDD  pch W=7.18u    L=0.24U
M3  QN  SIN   VSS      VSS    nch W=1.8u     L=0.24U
M4  VSS     Q   QN   VSS    nch W=1.8u     L=0.24U
M5  VDD  RIN    TP1    VDD  pch W=7.18u    L=0.24U
M6  TP1  QN   Q    VDD  pch W=7.18u    L=0.24U
M7  Q  QN   VSS      VSS    nch W=1.8u     L=0.24U
M8  VSS    RIN    Q    VSS    nch W=1.8u     L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lscs1 CLK DIN SETB CLRB QN Q
M18 Q TP5 VSS VSS nch W=1.88U L=0.24U
M11 TP5 TP4 TP2 VDD pch W=1.8U L=0.24U
M12 TP2 CLK TP5 VSS nch W=1.3U L=0.24U
M16 TP6 Q VSS VSS nch W=0.8U L=0.24U
M19 QN Q VDD VDD pch W=2.96U L=0.24U
M20 QN Q VSS VSS nch W=1.32U L=0.24U
M17 Q TP5 VDD VDD pch W=2.98U L=0.24U
M15 TP6 Q VDD VDD pch W=1.3U L=0.24U
M13 TP5 TP4 TP6 VSS nch W=0.8U L=0.24U
M14 TP6 CLK TP5 VDD pch W=1.8U L=0.24U
M9 TP4 CLK VDD VDD pch W=1.3U L=0.24U
M10 TP4 CLK VSS VSS nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 SETB VSS VSS nch W=0.8U L=0.24U
M5 TP2 CLRB VDD VDD pch W=2U L=0.24U
M4 TP2 DIN TP1 VDD pch W=2U L=0.24U
M6 TP2 CLRB TP3 VSS nch W=1U L=0.24U
M7 TP3 DIN VSS VSS nch W=1U L=0.24U
M8 TP3 TP0 VSS VSS nch W=1U L=0.24U
M3 TP1 TP0 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lscs2 CLK DIN SETB CLRB QN Q
M18 Q TP5 VSS VSS nch W=3.98U L=0.24U
M11 TP5 TP4 TP2 VDD pch W=2.8U L=0.24U
M12 TP2 CLK TP5 VSS nch W=2.6U L=0.24U
M16 TP6 Q VSS VSS nch W=0.8U L=0.24U
M19 QN Q VDD VDD pch W=5.96U L=0.24U
M20 QN Q VSS VSS nch W=2.42U L=0.24U
M17 Q TP5 VDD VDD pch W=6.02U L=0.24U
M15 TP6 Q VDD VDD pch W=1.3U L=0.24U
M13 TP5 TP4 TP6 VSS nch W=0.8U L=0.24U
M14 TP6 CLK TP5 VDD pch W=1.3U L=0.24U
M9 TP4 CLK VDD VDD pch W=1.3U L=0.24U
M10 TP4 CLK VSS VSS nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 SETB VSS VSS nch W=0.8U L=0.24U
M5 TP2 CLRB VDD VDD pch W=2.5U L=0.24U
M4 TP2 DIN TP1 VDD pch W=2.5U L=0.24U
M6 TP2 CLRB TP3 VSS nch W=1.3U L=0.24U
M7 TP3 DIN VSS VSS nch W=1.3U L=0.24U
M8 TP3 TP0 VSS VSS nch W=1.3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lss1 SETB DIN CLK QN Q
M11 Q TP2 VDD VDD pch W=3.14U L=0.24U
M12 Q SETB VDD VDD pch W=3.14U L=0.24U
M14 TP4 SETB VSS VSS nch W=2.88U L=0.24U
M13 Q TP2 TP4 VSS nch W=2.88U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M4 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M6 TP2 TP1 TP0 VDD pch W=2.2U L=0.24U
M5 TP0 CLK TP2 VSS nch W=1.8U L=0.24U
M8 TP2 TP1 TP3 VSS nch W=0.8U L=0.24U
M7 TP3 CLK TP2 VDD pch W=1.3U L=0.24U
M9 TP3 Q VDD VDD pch W=1.3U L=0.24U
M10 TP3 Q VSS VSS nch W=0.8U L=0.24U
M15 QN Q VDD VDD pch W=3.12U L=0.24U
M16 QN Q VSS VSS nch W=1.4U L=0.24U
M2 TP0 DIN VSS VSS nch W=0.9U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT lss2 SETB DIN CLK QN Q
M11 Q TP2 VDD VDD pch W=6.9U L=0.24U
M12 Q SETB VDD VDD pch W=6.9U L=0.24U
M14 TP4 SETB VSS VSS nch W=6.6U L=0.24U
M13 Q TP2 TP4 VSS nch W=6.6U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M4 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M6 TP2 TP1 TP0 VDD pch W=2.8U L=0.24U
M5 TP0 CLK TP2 VSS nch W=2.5U L=0.24U
M8 TP2 TP1 TP3 VSS nch W=0.8U L=0.24U
M7 TP3 CLK TP2 VDD pch W=1.3U L=0.24U
M9 TP3 Q VDD VDD pch W=1.3U L=0.24U
M10 TP3 Q VSS VSS nch W=0.8U L=0.24U
M15 QN Q VDD VDD pch W=6.8U L=0.24U
M16 QN Q VSS VSS nch W=3U L=0.24U
M2 TP0 DIN VSS VSS nch W=1.42U L=0.24U
M1 TP0 DIN VDD VDD pch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mx21s1 Q DIN1 SIN DIN2
M4 DIN2 SIN N1N438 VSS nch W=0.6U L=0.24U
M3 N1N438 N1N434 DIN1 VSS nch W=0.6U L=0.24U
M2 N1N434 SIN VSS VSS nch W=0.6U L=0.24U
M1 N1N434 SIN VDD VDD pch W=1.2U L=0.24U
M7 N1N441 N1N438 VSS VSS nch W=1U L=0.24U
M9 Q N1N441 VSS VSS nch W=1U L=0.24U
M6 N1N441 N1N438 VDD VDD pch W=1.3U L=0.24U
M8 Q N1N441 VDD VDD pch W=2.4U L=0.24U
M5 N1N438 N1N441 VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mux Q DIN1 SIN DIN2
M4 DIN2 SIN N1N438 VSS nch W=0.6U L=0.24U
M3 N1N438 N1N434 DIN1 VSS nch W=0.6U L=0.24U
M2 N1N434 SIN VSS VSS nch W=0.6U L=0.24U
M1 N1N434 SIN VDD VDD pch W=1.2U L=0.24U
M7 N1N441 N1N438 VSS VSS nch W=1U L=0.24U
M9 Q N1N441 VSS VSS nch W=1U L=0.24U
M6 N1N441 N1N438 VDD VDD pch W=1.3U L=0.24U
M8 Q N1N441 VDD VDD pch W=2.4U L=0.24U
M5 N1N438 N1N441 VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mx21s2 Q DIN1 SIN DIN2
M4 DIN2 SIN N1N438 VSS nch W=0.6U L=0.24U
M3 N1N438 N1N430 DIN2 VDD pch W=1.1U L=0.24U
M7 N1N498 N1N438 VDD VDD pch W=1.6U L=0.24U
M8 N1N498 N1N438 VSS VSS nch W=0.7U L=0.24U
M2 DIN1 N1N430 N1N438 VSS nch W=0.6U L=0.24U
M1 N1N438 SIN DIN1 VDD pch W=1.1U L=0.24U
M6 N1N430 SIN VSS VSS nch W=0.7U L=0.24U
M5 N1N430 SIN VDD VDD pch W=1.4U L=0.24U
M9 Q N1N498 VDD VDD pch W=3U L=0.24U
M10 Q N1N498 VSS VSS nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mx21s3 Q DIN1 SIN DIN2
M6 N1N430 SIN VSS VSS nch W=0.9U L=0.24U
M5 N1N430 SIN VDD VDD pch W=1.8U L=0.24U
M3 N1N438 N1N430 DIN2 VDD pch W=1.8U L=0.24U
M4 DIN2 SIN N1N438 VSS nch W=0.9U L=0.24U
M2 DIN1 N1N430 N1N438 VSS nch W=0.9U L=0.24U
M1 N1N438 SIN DIN1 VDD pch W=1.8U L=0.24U
M8 N1N483 N1N438 VSS VSS nch W=0.9U L=0.24U
M10 Q N1N483 VSS VSS nch W=3.6U L=0.24U
M7 N1N483 N1N438 VDD VDD pch W=2.2U L=0.24U
M9 Q N1N483 VDD VDD pch W=5.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mx41s1 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M3 N1N440 N1N429 DIN1 VSS nch W=0.8U L=0.24U
M4 N1N440 SIN0 DIN2 VSS nch W=0.8U L=0.24U
M5 N1N442 N1N429 DIN3 VSS nch W=0.8U L=0.24U
M6 N1N442 SIN0 DIN4 VSS nch W=0.8U L=0.24U
M10 N1N448 SIN1 N1N442 VSS nch W=0.6U L=0.24U
M9 N1N448 N1N451 N1N440 VSS nch W=0.6U L=0.24U
M2 N1N429 SIN0 VSS VSS nch W=0.6U L=0.24U
M1 N1N429 SIN0 VDD VDD pch W=1.2U L=0.24U
M7 N1N451 SIN1 VDD VDD pch W=1.2U L=0.24U
M8 N1N451 SIN1 VSS VSS nch W=0.6U L=0.24U
M13 N1N458 N1N448 VSS VSS nch W=1.1U L=0.24U
M12 N1N458 N1N448 VDD VDD pch W=2U L=0.24U
M14 Q N1N458 VDD VDD pch W=2.5U L=0.24U
M15 Q N1N458 VSS VSS nch W=1.3U L=0.24U
M11 N1N448 N1N458 VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mx41s2 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M2 DIN1 N1N564 N1N488 VSS nch W=0.8U L=0.24U
M1 N1N488 SIN0 DIN1 VDD pch W=1.6U L=0.24U
M3 N1N488 N1N564 DIN2 VDD pch W=1.6U L=0.24U
M4 DIN2 SIN0 N1N488 VSS nch W=0.8U L=0.24U
M5 N1N490 SIN0 DIN3 VDD pch W=1.6U L=0.24U
M6 DIN3 N1N564 N1N490 VSS nch W=0.8U L=0.24U
M7 N1N490 N1N564 DIN4 VDD pch W=1.6U L=0.24U
M8 DIN4 SIN0 N1N490 VSS nch W=0.8U L=0.24U
M10 N1N564 SIN0 VSS VSS nch W=0.8U L=0.24U
M9 N1N564 SIN0 VDD VDD pch W=1.6U L=0.24U
M11 N1N507 SIN1 VDD VDD pch W=1.2U L=0.24U
M12 N1N507 SIN1 VSS VSS nch W=0.6U L=0.24U
M15 N1N510 N1N507 N1N490 VDD pch W=1.2U L=0.24U
M16 N1N490 SIN1 N1N510 VSS nch W=0.6U L=0.24U
M13 N1N510 SIN1 N1N488 VDD pch W=1.2U L=0.24U
M14 N1N488 N1N507 N1N510 VSS nch W=0.6U L=0.24U
M17 N1N646 N1N510 VDD VDD pch W=2.4U L=0.24U
M19 Q N1N646 VDD VDD pch W=3.3U L=0.24U
M18 N1N646 N1N510 VSS VSS nch W=1U L=0.24U
M20 Q N1N646 VSS VSS nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mx41s3 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M14 N1N490 SIN1 N1N510 VSS nch W=0.9U L=0.24U
M13 N1N510 N1N507 N1N490 VDD pch W=1.8U L=0.24U
M2 DIN1 N1N493 N1N488 VSS nch W=1.2U L=0.24U
M1 N1N488 SIN0 DIN1 VDD pch W=2.4U L=0.24U
M4 DIN2 SIN0 N1N488 VSS nch W=1.2U L=0.24U
M3 N1N488 N1N493 DIN2 VDD pch W=2.4U L=0.24U
M5 N1N490 SIN0 DIN3 VDD pch W=2.4U L=0.24U
M6 DIN3 N1N493 N1N490 VSS nch W=1.2U L=0.24U
M7 N1N490 N1N493 DIN4 VDD pch W=2.4U L=0.24U
M8 DIN4 SIN0 N1N490 VSS nch W=1.2U L=0.24U
M11 N1N510 SIN1 N1N488 VDD pch W=1.8U L=0.24U
M12 N1N488 N1N507 N1N510 VSS nch W=0.9U L=0.24U
M17 Q N1N569 VDD VDD pch W=6.6U L=0.24U
M18 Q N1N569 VSS VSS nch W=4U L=0.24U
M10 N1N493 SIN0 VSS VSS nch W=1.2U L=0.24U
M9 N1N493 SIN0 VDD VDD pch W=2.5U L=0.24U
M19 N1N507 SIN1 VDD VDD pch W=1.8U L=0.24U
M20 N1N507 SIN1 VSS VSS nch W=0.9U L=0.24U
M15 N1N569 N1N510 VDD VDD pch W=3.5U L=0.24U
M16 N1N569 N1N510 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mxi21s1 Q DIN1 SIN DIN2
M4 DIN2 SIN N1N438 VSS nch W=0.6U L=0.24U
M7 Q N1N438 VSS VSS nch W=2.4U L=0.24U
M6 Q N1N438 VDD VDD pch W=2.4U L=0.24U
M1 N1N434 SIN VDD VDD pch W=1.2U L=0.24U
M2 N1N434 SIN VSS VSS nch W=0.6U L=0.24U
M3 N1N438 N1N434 DIN1 VSS nch W=0.6U L=0.24U
M5 N1N438 Q VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mxi21s2 Q DIN1 SIN DIN2
M8 Q N1N438 VSS VSS nch W=1.24U L=0.24U
M6 DIN2 SIN N1N438 VSS nch W=0.6U L=0.24U
M7 Q N1N438 VDD VDD pch W=3U L=0.24U
M5 N1N438 N1N430 DIN2 VDD pch W=1.1U L=0.24U
M4 DIN1 N1N430 N1N438 VSS nch W=0.6U L=0.24U
M3 N1N438 SIN DIN1 VDD pch W=1.1U L=0.24U
M2 N1N430 SIN VSS VSS nch W=0.7U L=0.24U
M1 N1N430 SIN VDD VDD pch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mxi21s3 Q DIN1 SIN DIN2
M8 Q N1N438 VSS VSS nch W=2.1U L=0.24U
M6 DIN2 SIN N1N438 VSS nch W=0.9U L=0.24U
M7 Q N1N438 VDD VDD pch W=5.7U L=0.24U
M5 N1N438 N1N430 DIN2 VDD pch W=1.8U L=0.24U
M4 DIN1 N1N430 N1N438 VSS nch W=0.9U L=0.24U
M3 N1N438 SIN DIN1 VDD pch W=1.8U L=0.24U
M2 N1N430 SIN VSS VSS nch W=0.9U L=0.24U
M1 N1N430 SIN VDD VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mxi41s1 Q DIN1 SIN0 SIN1 DIN2 DIN3 DIN4
M3 N1N440 N1N429 DIN1 VSS nch W=0.8U L=0.24U
M4 N1N440 SIN0 DIN2 VSS nch W=0.8U L=0.24U
M5 N1N442 N1N429 DIN3 VSS nch W=0.8U L=0.24U
M6 N1N442 SIN0 DIN4 VSS nch W=0.8U L=0.24U
M10 N1N448 SIN1 N1N442 VSS nch W=0.6U L=0.24U
M9 N1N448 N1N451 N1N440 VSS nch W=0.6U L=0.24U
M13 Q N1N448 VSS VSS nch W=1.7U L=0.24U
M12 Q N1N448 VDD VDD pch W=2.5U L=0.24U
M2 N1N429 SIN0 VSS VSS nch W=0.6U L=0.24U
M1 N1N429 SIN0 VDD VDD pch W=1.2U L=0.24U
M8 N1N451 SIN1 VSS VSS nch W=0.6U L=0.24U
M7 N1N451 SIN1 VDD VDD pch W=1.2U L=0.24U
M11 N1N448 Q VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mxi41s2 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M18 Q N1N510 VSS VSS nch W=1.5U L=0.24U
M16 N1N490 SIN1 N1N510 VSS nch W=0.6U L=0.24U
M15 N1N510 N1N589 N1N490 VDD pch W=1.2U L=0.24U
M17 Q N1N510 VDD VDD pch W=3.4U L=0.24U
M2 DIN1 N1N493 N1N488 VSS nch W=0.8U L=0.24U
M1 N1N488 SIN0 DIN1 VDD pch W=1.6U L=0.24U
M4 DIN2 SIN0 N1N488 VSS nch W=0.8U L=0.24U
M3 N1N488 N1N493 DIN2 VDD pch W=1.6U L=0.24U
M6 DIN3 N1N493 N1N490 VSS nch W=0.8U L=0.24U
M5 N1N490 SIN0 DIN3 VDD pch W=1.6U L=0.24U
M8 DIN4 SIN0 N1N490 VSS nch W=0.8U L=0.24U
M7 N1N490 N1N493 DIN4 VDD pch W=1.6U L=0.24U
M9 N1N493 SIN0 VDD VDD pch W=1.6U L=0.24U
M10 N1N493 SIN0 VSS VSS nch W=0.8U L=0.24U
M11 N1N589 SIN1 VDD VDD pch W=1.2U L=0.24U
M12 N1N589 SIN1 VSS VSS nch W=0.6U L=0.24U
M14 N1N488 N1N589 N1N510 VSS nch W=0.6U L=0.24U
M13 N1N510 SIN1 N1N488 VDD pch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT mxi41s3 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M18 Q N1N510 VSS VSS nch W=2.2U L=0.24U
M16 N1N490 SIN1 N1N510 VSS nch W=0.9U L=0.24U
M15 N1N510 N1N589 N1N490 VDD pch W=1.8U L=0.24U
M17 Q N1N510 VDD VDD pch W=5.7U L=0.24U
M2 DIN1 N1N493 N1N488 VSS nch W=1.2U L=0.24U
M1 N1N488 SIN0 DIN1 VDD pch W=2.4U L=0.24U
M4 DIN2 SIN0 N1N488 VSS nch W=1.2U L=0.24U
M3 N1N488 N1N493 DIN2 VDD pch W=2.4U L=0.24U
M6 DIN3 N1N493 N1N490 VSS nch W=1.2U L=0.24U
M5 N1N490 SIN0 DIN3 VDD pch W=2.4U L=0.24U
M8 DIN4 SIN0 N1N490 VSS nch W=1.2U L=0.24U
M7 N1N490 N1N493 DIN4 VDD pch W=2.4U L=0.24U
M9 N1N493 SIN0 VDD VDD pch W=2.5U L=0.24U
M10 N1N493 SIN0 VSS VSS nch W=1.2U L=0.24U
M11 N1N589 SIN1 VDD VDD pch W=1.8U L=0.24U
M12 N1N589 SIN1 VSS VSS nch W=0.9U L=0.24U
M14 N1N488 N1N589 N1N510 VSS nch W=0.9U L=0.24U
M13 N1N510 SIN1 N1N488 VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s1 Q DIN
M4 Q N1N262 VSS VSS nch W=1.5U L=0.24U
M3 Q N1N262 VDD VDD pch W=2.5U L=0.24U
M1 N1N262 DIN VDD VDD pch W=2.1U L=0.24U
M2 N1N262 DIN VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s10 Q DIN
M4 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M3 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M1 N1N318 DIN VDD VDD pch W=43U L=0.24U
M2 N1N318 DIN VSS VSS nch W=20U L=0.24U
M6 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M5 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M7 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M8 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M10 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M9 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M11 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M12 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M14 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M13 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M15 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M16 Q N1N318 VSS VSS nch W=3.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s11 DIN Q
M4 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M3 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M1 N1N318 DIN VDD VDD pch W=53U L=0.24U
M2 N1N318 DIN VSS VSS nch W=24U L=0.24U
M6 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M5 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M7 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M8 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M10 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M9 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M11 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M12 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M14 Q N1N318 VSS VSS nch W=3.5U L=0.24U
M13 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M15 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M16 Q N1N318 VSS VSS nch W=3.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s12 DIN Q
M4 Q N1N318 VSS VSS nch W=3.7U L=0.24U
M3 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M1 N1N318 DIN VDD VDD pch W=55U L=0.24U
M2 N1N318 DIN VSS VSS nch W=27U L=0.24U
M6 Q N1N318 VSS VSS nch W=3.7U L=0.24U
M5 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M7 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M8 Q N1N318 VSS VSS nch W=3.7U L=0.24U
M10 Q N1N318 VSS VSS nch W=3.7U L=0.24U
M9 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M11 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M12 Q N1N318 VSS VSS nch W=3.7U L=0.24U
M14 Q N1N318 VSS VSS nch W=3.7U L=0.24U
M13 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M15 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M16 Q N1N318 VSS VSS nch W=3.7U L=0.24U
M17 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M18 Q N1N318 VSS VSS nch W=3.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s2 Q DIN
M4 Q N1N262 VSS VSS nch W=1.5U L=0.24U
M3 Q N1N262 VDD VDD pch W=2.8U L=0.24U
M1 N1N262 DIN VDD VDD pch W=2.5U L=0.24U
M2 N1N262 DIN VSS VSS nch W=1.4U L=0.24U
M6 Q N1N262 VSS VSS nch W=1.5U L=0.24U
M5 Q N1N262 VDD VDD pch W=2.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s3 Q DIN
M4 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M3 Q N1N262 VDD VDD pch W=2.3U L=0.24U
M1 N1N262 DIN VDD VDD pch W=3.9U L=0.24U
M2 N1N262 DIN VSS VSS nch W=1.6U L=0.24U
M6 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M5 Q N1N262 VDD VDD pch W=2.3U L=0.24U
M7 Q N1N262 VDD VDD pch W=2.3U L=0.24U
M8 Q N1N262 VSS VSS nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s4 Q DIN
M4 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M3 Q N1N262 VDD VDD pch W=2U L=0.24U
M1 N1N262 DIN VDD VDD pch W=4U L=0.24U
M2 N1N262 DIN VSS VSS nch W=2U L=0.24U
M6 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M5 Q N1N262 VDD VDD pch W=2U L=0.24U
M7 Q N1N262 VDD VDD pch W=2U L=0.24U
M8 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M10 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M9 Q N1N262 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s5 Q DIN
M4 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M3 Q N1N262 VDD VDD pch W=2U L=0.24U
M1 N1N262 DIN VDD VDD pch W=5.5U L=0.24U
M2 N1N262 DIN VSS VSS nch W=2.6U L=0.24U
M6 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M5 Q N1N262 VDD VDD pch W=2U L=0.24U
M7 Q N1N262 VDD VDD pch W=2U L=0.24U
M8 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M10 Q N1N262 VSS VSS nch W=1.1U L=0.24U
M9 Q N1N262 VDD VDD pch W=2U L=0.24U
M11 Q N1N262 VDD VDD pch W=2U L=0.24U
M12 Q N1N262 VSS VSS nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s6 Q DIN
M4 Q N1N318 VSS VSS nch W=1.1U L=0.24U
M3 Q N1N318 VDD VDD pch W=2U L=0.24U
M1 N1N318 DIN VDD VDD pch W=6.2U L=0.24U
M2 N1N318 DIN VSS VSS nch W=3U L=0.24U
M6 Q N1N318 VSS VSS nch W=1.1U L=0.24U
M5 Q N1N318 VDD VDD pch W=2U L=0.24U
M7 Q N1N318 VDD VDD pch W=2U L=0.24U
M8 Q N1N318 VSS VSS nch W=1.1U L=0.24U
M10 Q N1N318 VSS VSS nch W=1.1U L=0.24U
M9 Q N1N318 VDD VDD pch W=2U L=0.24U
M11 Q N1N318 VDD VDD pch W=2U L=0.24U
M12 Q N1N318 VSS VSS nch W=1.1U L=0.24U
M14 Q N1N318 VSS VSS nch W=1.1U L=0.24U
M13 Q N1N318 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s7 DIN Q
M4 Q N1N318 VSS VSS nch W=1.7U L=0.24U
M3 Q N1N318 VDD VDD pch W=3U L=0.24U
M1 N1N318 DIN VDD VDD pch W=8U L=0.24U
M2 N1N318 DIN VSS VSS nch W=3.8U L=0.24U
M6 Q N1N318 VSS VSS nch W=1.7U L=0.24U
M5 Q N1N318 VDD VDD pch W=3U L=0.24U
M7 Q N1N318 VDD VDD pch W=3U L=0.24U
M8 Q N1N318 VSS VSS nch W=1.7U L=0.24U
M10 Q N1N318 VSS VSS nch W=1.7U L=0.24U
M9 Q N1N318 VDD VDD pch W=3U L=0.24U
M11 Q N1N318 VDD VDD pch W=3U L=0.24U
M12 Q N1N318 VSS VSS nch W=1.7U L=0.24U
M14 Q N1N318 VSS VSS nch W=1.7U L=0.24U
M13 Q N1N318 VDD VDD pch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s8 DIN Q
M4 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M3 Q N1N318 VDD VDD pch W=4U L=0.24U
M1 N1N318 DIN VDD VDD pch W=15U L=0.24U
M2 N1N318 DIN VSS VSS nch W=7U L=0.24U
M6 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M5 Q N1N318 VDD VDD pch W=4U L=0.24U
M7 Q N1N318 VDD VDD pch W=4U L=0.24U
M8 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M10 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M9 Q N1N318 VDD VDD pch W=4U L=0.24U
M11 Q N1N318 VDD VDD pch W=4U L=0.24U
M12 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M14 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M13 Q N1N318 VDD VDD pch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nb1s9 DIN Q
M4 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M3 Q N1N318 VDD VDD pch W=4U L=0.24U
M1 N1N318 DIN VDD VDD pch W=26U L=0.24U
M2 N1N318 DIN VSS VSS nch W=12U L=0.24U
M6 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M5 Q N1N318 VDD VDD pch W=4U L=0.24U
M7 Q N1N318 VDD VDD pch W=4U L=0.24U
M8 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M10 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M9 Q N1N318 VDD VDD pch W=4U L=0.24U
M11 Q N1N318 VDD VDD pch W=4U L=0.24U
M12 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M14 Q N1N318 VSS VSS nch W=2.3U L=0.24U
M13 Q N1N318 VDD VDD pch W=4U L=0.24U
M15 Q N1N318 VDD VDD pch W=4U L=0.24U
M16 Q N1N318 VSS VSS nch W=2.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd2s1 Q DIN1 DIN2
M3 Q DIN1 N1N275 VSS nch W=1.16U L=0.24U
M1 Q DIN1 VDD VDD pch W=1.8U L=0.24U
M2 VDD DIN2 Q VDD pch W=1.8U L=0.24U
M4 N1N275 DIN2 VSS VSS nch W=1.16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd2s2 Q DIN1 DIN2
M3 Q DIN1 N1N275 VSS nch W=2.18U L=0.24U
M1 Q DIN1 VDD VDD pch W=3.3U L=0.24U
M2 VDD DIN2 Q VDD pch W=3.3U L=0.24U
M4 N1N275 DIN2 VSS VSS nch W=2.18U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd2s3 Q DIN1 DIN2
M3 Q DIN1 N1N275 VSS nch W=4U L=0.24U
M1 Q DIN1 VDD VDD pch W=5.9U L=0.24U
M2 VDD DIN2 Q VDD pch W=5.9U L=0.24U
M4 N1N275 DIN2 VSS VSS nch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd3s1 Q DIN1 DIN2 DIN3
M4 Q DIN1 N1N260 VSS nch W=1.5U L=0.24U
M3 Q DIN3 VDD VDD pch W=1.8U L=0.24U
M2 Q DIN2 VDD VDD pch W=1.8U L=0.24U
M1 Q DIN1 VDD VDD pch W=1.8U L=0.24U
M6 N1N293 DIN3 VSS VSS nch W=1.5U L=0.24U
M5 N1N260 DIN2 N1N293 VSS nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd3s2 Q DIN1 DIN2 DIN3
M4 Q DIN1 N1N260 VSS nch W=2.64U L=0.24U
M3 Q DIN3 VDD VDD pch W=3.12U L=0.24U
M2 Q DIN2 VDD VDD pch W=3.12U L=0.24U
M1 Q DIN1 VDD VDD pch W=3.12U L=0.24U
M6 N1N293 DIN3 VSS VSS nch W=2.64U L=0.24U
M5 N1N260 DIN2 N1N293 VSS nch W=2.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd3s3 Q DIN1 DIN2 DIN3
M4 Q DIN1 N1N260 VSS nch W=4.8U L=0.24U
M3 Q DIN3 VDD VDD pch W=6U L=0.24U
M2 Q DIN2 VDD VDD pch W=6U L=0.24U
M1 Q DIN1 VDD VDD pch W=6U L=0.24U
M6 N1N293 DIN3 VSS VSS nch W=5.6U L=0.24U
M5 N1N260 DIN2 N1N293 VSS nch W=5.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd4s1 Q DIN1 DIN2 DIN3 DIN4
M1 Q DIN1 VDD VDD pch W=1.9U L=0.24U
M2 Q DIN2 VDD VDD pch W=1.9U L=0.24U
M3 Q DIN3 VDD VDD pch W=1.9U L=0.24U
M4 Q DIN4 VDD VDD pch W=1.9U L=0.24U
M5 Q DIN1 N1N348 VSS nch W=1.8U L=0.24U
M6 N1N348 DIN2 N1N347 VSS nch W=1.84U L=0.24U
M7 N1N347 DIN3 N1N346 VSS nch W=1.94U L=0.24U
M8 N1N346 DIN4 VSS VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd4s2 Q DIN1 DIN2 DIN3 DIN4
M1 Q DIN1 VDD VDD pch W=3.12U L=0.24U
M2 Q DIN2 VDD VDD pch W=3.12U L=0.24U
M3 Q DIN3 VDD VDD pch W=3.12U L=0.24U
M4 Q DIN4 VDD VDD pch W=3.12U L=0.24U
M5 Q DIN1 N1N348 VSS nch W=2.98U L=0.24U
M6 N1N348 DIN2 N1N347 VSS nch W=3U L=0.24U
M7 N1N347 DIN3 N1N346 VSS nch W=3.1U L=0.24U
M8 N1N346 DIN4 VSS VSS nch W=3.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nnd4s3 Q DIN1 DIN2 DIN3 DIN4
M4 N1N280 DIN2 VSS VSS nch W=4.1U L=0.24U
M3 N1N269 DIN1 N1N280 VSS nch W=3.1U L=0.24U
M14 Q N1N315 VSS VSS nch W=4U L=0.24U
M12 VSS N1N298 N1N315 VSS nch W=3.1U L=0.24U
M11 N1N315 N1N269 VSS VSS nch W=3.1U L=0.24U
M8 N1N309 DIN4 VSS VSS nch W=4.1U L=0.24U
M7 N1N298 DIN3 N1N309 VSS nch W=3.1U L=0.24U
M5 N1N298 DIN3 VDD VDD pch W=3.7U L=0.24U
M6 VDD DIN4 N1N298 VDD pch W=3.7U L=0.24U
M10 N1N325 N1N298 N1N315 VDD pch W=7.2U L=0.24U
M1 N1N269 DIN1 VDD VDD pch W=3.7U L=0.24U
M2 VDD DIN2 N1N269 VDD pch W=3.7U L=0.24U
M9 N1N325 N1N269 VDD VDD pch W=7.5U L=0.24U
M13 Q N1N315 VDD VDD pch W=8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and5s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M4 N1N442 DIN1 N1N438 VSS nch W=3.9U L=0.24U
M1 N1N442 DIN1 VDD VDD pch W=4.2U L=0.24U
M2 N1N442 DIN2 VDD VDD pch W=4.2U L=0.24U
M3 N1N442 DIN3 VDD VDD pch W=4.2U L=0.24U
M5 N1N438 DIN2 N1N440 VSS nch W=4.8U L=0.24U
M6 N1N440 DIN3 VSS VSS nch W=5.8U L=0.24U
M11 N1N446 N1N442 VDD VDD pch W=6.7U L=0.24U
M12 N1N446 N1N455 N1N448 VDD pch W=6.1U L=0.24U
M13 N1N448 N1N442 VSS VSS nch W=3.1U L=0.24U
M14 VSS N1N455 N1N448 VSS nch W=3.1U L=0.24U
M7 N1N455 DIN4 VDD VDD pch W=4.2U L=0.24U
M8 N1N455 DIN5 VDD VDD pch W=4.2U L=0.24U
M9 N1N455 DIN4 N1N457 VSS nch W=3.4U L=0.24U
M10 N1N457 DIN5 VSS VSS nch W=3.9U L=0.24U
M15 Q N1N448 VDD VDD pch W=4.3U L=0.24U
M16 Q N1N448 VSS VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nnd5s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M4 N1N442 DIN1 N1N438 VSS nch W=3.9U L=0.24U
M1 N1N442 DIN1 VDD VDD pch W=4.2U L=0.24U
M2 N1N442 DIN2 VDD VDD pch W=4.2U L=0.24U
M3 N1N442 DIN3 VDD VDD pch W=4.2U L=0.24U
M5 N1N438 DIN2 N1N440 VSS nch W=4.8U L=0.24U
M6 N1N440 DIN3 VSS VSS nch W=5.8U L=0.24U
M11 N1N446 N1N442 VDD VDD pch W=6.7U L=0.24U
M12 N1N446 N1N455 N1N448 VDD pch W=6.1U L=0.24U
M13 N1N448 N1N442 VSS VSS nch W=3.1U L=0.24U
M14 VSS N1N455 N1N448 VSS nch W=3.1U L=0.24U
M7 N1N455 DIN4 VDD VDD pch W=4.2U L=0.24U
M8 N1N455 DIN5 VDD VDD pch W=4.2U L=0.24U
M9 N1N455 DIN4 N1N457 VSS nch W=3.4U L=0.24U
M10 N1N457 DIN5 VSS VSS nch W=3.9U L=0.24U
M15 Q N1N448 VDD VDD pch W=4.3U L=0.24U
M16 Q N1N448 VSS VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nnd5s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M4 N1N442 DIN1 N1N438 VSS nch W=3.9U L=0.24U
M1 N1N442 DIN1 VDD VDD pch W=4.2U L=0.24U
M2 N1N442 DIN2 VDD VDD pch W=4.2U L=0.24U
M3 N1N442 DIN3 VDD VDD pch W=4.2U L=0.24U
M5 N1N438 DIN2 N1N440 VSS nch W=4.8U L=0.24U
M6 N1N440 DIN3 VSS VSS nch W=5.8U L=0.24U
M11 N1N446 N1N442 VDD VDD pch W=6.7U L=0.24U
M12 N1N446 N1N455 N1N448 VDD pch W=6.1U L=0.24U
M13 N1N448 N1N442 VSS VSS nch W=3.1U L=0.24U
M14 VSS N1N455 N1N448 VSS nch W=3.1U L=0.24U
M7 N1N455 DIN4 VDD VDD pch W=4.2U L=0.24U
M8 N1N455 DIN5 VDD VDD pch W=4.2U L=0.24U
M9 N1N455 DIN4 N1N457 VSS nch W=3.4U L=0.24U
M10 N1N457 DIN5 VSS VSS nch W=3.9U L=0.24U
M15 Q N1N448 VDD VDD pch W=4.3U L=0.24U
M16 Q N1N448 VSS VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and6s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M1 N1N419 DIN1 VDD VDD pch W=4.1U L=0.24U
M2 N1N419 DIN2 VDD VDD pch W=4.1U L=0.24U
M3 N1N419 DIN3 VDD VDD pch W=4.1U L=0.24U
M4 N1N419 DIN1 N1N429 VSS nch W=3.9U L=0.24U
M5 N1N429 DIN2 N1N428 VSS nch W=4.8U L=0.24U
M6 N1N428 DIN3 VSS VSS nch W=5.8U L=0.24U
M13 N1N427 N1N419 VDD VDD pch W=6.7U L=0.24U
M14 N1N427 N1N424 N1N425 VDD pch W=6.1U L=0.24U
M15 N1N425 N1N419 VSS VSS nch W=3U L=0.24U
M16 VSS N1N424 N1N425 VSS nch W=3U L=0.24U
M10 N1N424 DIN4 N1N453 VSS nch W=3.9U L=0.24U
M7 N1N424 DIN4 VDD VDD pch W=4.1U L=0.24U
M8 N1N424 DIN5 VDD VDD pch W=4.1U L=0.24U
M9 N1N424 DIN6 VDD VDD pch W=4.1U L=0.24U
M11 N1N453 DIN5 N1N455 VSS nch W=4.8U L=0.24U
M12 N1N455 DIN6 VSS VSS nch W=5.8U L=0.24U
M18 Q N1N425 VSS VSS nch W=2.1U L=0.24U
M17 Q N1N425 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nnd6s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M1 N1N419 DIN1 VDD VDD pch W=4.1U L=0.24U
M2 N1N419 DIN2 VDD VDD pch W=4.1U L=0.24U
M3 N1N419 DIN3 VDD VDD pch W=4.1U L=0.24U
M4 N1N419 DIN1 N1N429 VSS nch W=3.9U L=0.24U
M5 N1N429 DIN2 N1N428 VSS nch W=4.8U L=0.24U
M6 N1N428 DIN3 VSS VSS nch W=5.8U L=0.24U
M13 N1N427 N1N419 VDD VDD pch W=6.7U L=0.24U
M14 N1N427 N1N424 N1N425 VDD pch W=6.1U L=0.24U
M15 N1N425 N1N419 VSS VSS nch W=3U L=0.24U
M16 VSS N1N424 N1N425 VSS nch W=3U L=0.24U
M10 N1N424 DIN4 N1N453 VSS nch W=3.9U L=0.24U
M7 N1N424 DIN4 VDD VDD pch W=4.1U L=0.24U
M8 N1N424 DIN5 VDD VDD pch W=4.1U L=0.24U
M9 N1N424 DIN6 VDD VDD pch W=4.1U L=0.24U
M11 N1N453 DIN5 N1N455 VSS nch W=4.8U L=0.24U
M12 N1N455 DIN6 VSS VSS nch W=5.8U L=0.24U
M18 Q N1N425 VSS VSS nch W=2.1U L=0.24U
M17 Q N1N425 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and7s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M1 N1N439 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N439 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 VDD DIN3 N1N439 VDD pch W=2.1U L=0.24U
M4 N1N439 DIN1 N1N425 VSS nch W=2.4U L=0.24U
M5 N1N425 DIN2 N1N424 VSS nch W=2.6U L=0.24U
M6 N1N424 DIN3 VSS VSS nch W=2.8U L=0.24U
M11 N1N448 DIN7 VDD VDD pch W=2.1U L=0.24U
M12 N1N448 DIN6 VDD VDD pch W=2.1U L=0.24U
M13 VDD DIN5 N1N448 VDD pch W=2.1U L=0.24U
M14 VDD DIN4 N1N448 VDD pch W=2.1U L=0.24U
M15 N1N448 DIN4 N1N423 VSS nch W=6.3U L=0.24U
M16 N1N423 DIN5 N1N422 VSS nch W=6.5U L=0.24U
M17 N1N422 DIN6 N1N421 VSS nch W=6.7U L=0.24U
M18 N1N421 DIN7 VSS VSS nch W=6.9U L=0.24U
M7 N1N454 N1N439 VDD VDD pch W=5.2U L=0.24U
M8 N1N454 N1N448 N1N455 VDD pch W=5.2U L=0.24U
M9 N1N455 N1N439 VSS VSS nch W=2.3U L=0.24U
M10 VSS N1N448 N1N455 VSS nch W=2.3U L=0.24U
M20 Q N1N455 VSS VSS nch W=2.4U L=0.24U
M19 Q N1N455 VDD VDD pch W=6.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nnd7s3 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M1 N1N439 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N439 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 VDD DIN3 N1N439 VDD pch W=2.1U L=0.24U
M4 N1N439 DIN1 N1N425 VSS nch W=2.4U L=0.24U
M5 N1N425 DIN2 N1N424 VSS nch W=2.6U L=0.24U
M6 N1N424 DIN3 VSS VSS nch W=2.8U L=0.24U
M11 N1N448 DIN7 VDD VDD pch W=2.1U L=0.24U
M12 N1N448 DIN6 VDD VDD pch W=2.1U L=0.24U
M13 VDD DIN5 N1N448 VDD pch W=2.1U L=0.24U
M14 VDD DIN4 N1N448 VDD pch W=2.1U L=0.24U
M15 N1N448 DIN4 N1N423 VSS nch W=6.3U L=0.24U
M16 N1N423 DIN5 N1N422 VSS nch W=6.5U L=0.24U
M17 N1N422 DIN6 N1N421 VSS nch W=6.7U L=0.24U
M18 N1N421 DIN7 VSS VSS nch W=6.9U L=0.24U
M7 N1N454 N1N439 VDD VDD pch W=5.2U L=0.24U
M8 N1N454 N1N448 N1N455 VDD pch W=5.2U L=0.24U
M9 N1N455 N1N439 VSS VSS nch W=2.3U L=0.24U
M10 VSS N1N448 N1N455 VSS nch W=2.3U L=0.24U
M20 Q N1N455 VSS VSS nch W=2.4U L=0.24U
M19 Q N1N455 VDD VDD pch W=6.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or8s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 Q
M5 N1N304 DIN1 N1N314 VSS nch W=6.3U L=0.24U
M1 N1N304 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N304 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 N1N304 DIN3 VDD VDD pch W=2.1U L=0.24U
M4 N1N304 DIN4 VDD VDD pch W=2.1U L=0.24U
M6 N1N314 DIN2 N1N316 VSS nch W=6.5U L=0.24U
M7 N1N316 DIN3 N1N318 VSS nch W=6.7U L=0.24U
M8 N1N318 DIN4 VSS VSS nch W=6.9U L=0.24U
M9 N1N343 N1N304 VDD VDD pch W=5.4U L=0.24U
M10 N1N343 N1N413 N1N345 VDD pch W=5.4U L=0.24U
M11 N1N345 N1N304 VSS VSS nch W=1.5U L=0.24U
M12 VSS N1N413 N1N345 VSS nch W=1.5U L=0.24U
M13 N1N413 DIN5 VDD VDD pch W=2.1U L=0.24U
M14 N1N413 DIN6 VDD VDD pch W=2.1U L=0.24U
M15 N1N413 DIN7 VDD VDD pch W=2.1U L=0.24U
M16 N1N413 DIN8 VDD VDD pch W=2.1U L=0.24U
M17 N1N413 DIN5 N1N362 VSS nch W=6.3U L=0.24U
M18 N1N362 DIN6 N1N364 VSS nch W=6.5U L=0.24U
M19 N1N364 DIN7 N1N366 VSS nch W=6.7U L=0.24U
M20 N1N366 DIN8 VSS VSS nch W=6.9U L=0.24U
M22 Q N1N345 VSS VSS nch W=3U L=0.24U
M21 Q N1N345 VDD VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT xor8s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 Q
M5 N1N304 DIN1 N1N314 VSS nch W=6.3U L=0.24U
M1 N1N304 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N304 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 N1N304 DIN3 VDD VDD pch W=2.1U L=0.24U
M4 N1N304 DIN4 VDD VDD pch W=2.1U L=0.24U
M6 N1N314 DIN2 N1N316 VSS nch W=6.5U L=0.24U
M7 N1N316 DIN3 N1N318 VSS nch W=6.7U L=0.24U
M8 N1N318 DIN4 VSS VSS nch W=6.9U L=0.24U
M9 N1N343 N1N304 VDD VDD pch W=5.4U L=0.24U
M10 N1N343 N1N413 N1N345 VDD pch W=5.4U L=0.24U
M11 N1N345 N1N304 VSS VSS nch W=1.5U L=0.24U
M12 VSS N1N413 N1N345 VSS nch W=1.5U L=0.24U
M13 N1N413 DIN5 VDD VDD pch W=2.1U L=0.24U
M14 N1N413 DIN6 VDD VDD pch W=2.1U L=0.24U
M15 N1N413 DIN7 VDD VDD pch W=2.1U L=0.24U
M16 N1N413 DIN8 VDD VDD pch W=2.1U L=0.24U
M17 N1N413 DIN5 N1N362 VSS nch W=6.3U L=0.24U
M18 N1N362 DIN6 N1N364 VSS nch W=6.5U L=0.24U
M19 N1N364 DIN7 N1N366 VSS nch W=6.7U L=0.24U
M20 N1N366 DIN8 VSS VSS nch W=6.9U L=0.24U
M22 Q N1N345 VSS VSS nch W=3U L=0.24U
M21 Q N1N345 VDD VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT xnr8s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 Q
M5 N1N304 DIN1 N1N314 VSS nch W=6.3U L=0.24U
M1 N1N304 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N304 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 N1N304 DIN3 VDD VDD pch W=2.1U L=0.24U
M4 N1N304 DIN4 VDD VDD pch W=2.1U L=0.24U
M6 N1N314 DIN2 N1N316 VSS nch W=6.5U L=0.24U
M7 N1N316 DIN3 N1N318 VSS nch W=6.7U L=0.24U
M8 N1N318 DIN4 VSS VSS nch W=6.9U L=0.24U
M9 N1N343 N1N304 VDD VDD pch W=5.4U L=0.24U
M10 N1N343 N1N413 N1N345 VDD pch W=5.4U L=0.24U
M11 N1N345 N1N304 VSS VSS nch W=1.5U L=0.24U
M12 VSS N1N413 N1N345 VSS nch W=1.5U L=0.24U
M13 N1N413 DIN5 VDD VDD pch W=2.1U L=0.24U
M14 N1N413 DIN6 VDD VDD pch W=2.1U L=0.24U
M15 N1N413 DIN7 VDD VDD pch W=2.1U L=0.24U
M16 N1N413 DIN8 VDD VDD pch W=2.1U L=0.24U
M17 N1N413 DIN5 N1N362 VSS nch W=6.3U L=0.24U
M18 N1N362 DIN6 N1N364 VSS nch W=6.5U L=0.24U
M19 N1N364 DIN7 N1N366 VSS nch W=6.7U L=0.24U
M20 N1N366 DIN8 VSS VSS nch W=6.9U L=0.24U
M22 Q N1N345 VSS VSS nch W=3U L=0.24U
M21 Q N1N345 VDD VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nor8s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 Q
M5 N1N304 DIN1 N1N314 VSS nch W=6.3U L=0.24U
M1 N1N304 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N304 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 N1N304 DIN3 VDD VDD pch W=2.1U L=0.24U
M4 N1N304 DIN4 VDD VDD pch W=2.1U L=0.24U
M6 N1N314 DIN2 N1N316 VSS nch W=6.5U L=0.24U
M7 N1N316 DIN3 N1N318 VSS nch W=6.7U L=0.24U
M8 N1N318 DIN4 VSS VSS nch W=6.9U L=0.24U
M9 N1N343 N1N304 VDD VDD pch W=5.4U L=0.24U
M10 N1N343 N1N413 N1N345 VDD pch W=5.4U L=0.24U
M11 N1N345 N1N304 VSS VSS nch W=1.5U L=0.24U
M12 VSS N1N413 N1N345 VSS nch W=1.5U L=0.24U
M13 N1N413 DIN5 VDD VDD pch W=2.1U L=0.24U
M14 N1N413 DIN6 VDD VDD pch W=2.1U L=0.24U
M15 N1N413 DIN7 VDD VDD pch W=2.1U L=0.24U
M16 N1N413 DIN8 VDD VDD pch W=2.1U L=0.24U
M17 N1N413 DIN5 N1N362 VSS nch W=6.3U L=0.24U
M18 N1N362 DIN6 N1N364 VSS nch W=6.5U L=0.24U
M19 N1N364 DIN7 N1N366 VSS nch W=6.7U L=0.24U
M20 N1N366 DIN8 VSS VSS nch W=6.9U L=0.24U
M22 Q N1N345 VSS VSS nch W=3U L=0.24U
M21 Q N1N345 VDD VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nnd8s3 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 Q
M5 N1N304 DIN1 N1N314 VSS nch W=6.3U L=0.24U
M1 N1N304 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N304 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 N1N304 DIN3 VDD VDD pch W=2.1U L=0.24U
M4 N1N304 DIN4 VDD VDD pch W=2.1U L=0.24U
M6 N1N314 DIN2 N1N316 VSS nch W=6.5U L=0.24U
M7 N1N316 DIN3 N1N318 VSS nch W=6.7U L=0.24U
M8 N1N318 DIN4 VSS VSS nch W=6.9U L=0.24U
M9 N1N343 N1N304 VDD VDD pch W=5.4U L=0.24U
M10 N1N343 N1N413 N1N345 VDD pch W=5.4U L=0.24U
M11 N1N345 N1N304 VSS VSS nch W=1.5U L=0.24U
M12 VSS N1N413 N1N345 VSS nch W=1.5U L=0.24U
M13 N1N413 DIN5 VDD VDD pch W=2.1U L=0.24U
M14 N1N413 DIN6 VDD VDD pch W=2.1U L=0.24U
M15 N1N413 DIN7 VDD VDD pch W=2.1U L=0.24U
M16 N1N413 DIN8 VDD VDD pch W=2.1U L=0.24U
M17 N1N413 DIN5 N1N362 VSS nch W=6.3U L=0.24U
M18 N1N362 DIN6 N1N364 VSS nch W=6.5U L=0.24U
M19 N1N364 DIN7 N1N366 VSS nch W=6.7U L=0.24U
M20 N1N366 DIN8 VSS VSS nch W=6.9U L=0.24U
M22 Q N1N345 VSS VSS nch W=3U L=0.24U
M21 Q N1N345 VDD VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and8s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 Q
M5 N1N304 DIN1 N1N314 VSS nch W=6.3U L=0.24U
M1 N1N304 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N304 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 N1N304 DIN3 VDD VDD pch W=2.1U L=0.24U
M4 N1N304 DIN4 VDD VDD pch W=2.1U L=0.24U
M6 N1N314 DIN2 N1N316 VSS nch W=6.5U L=0.24U
M7 N1N316 DIN3 N1N318 VSS nch W=6.7U L=0.24U
M8 N1N318 DIN4 VSS VSS nch W=6.9U L=0.24U
M9 N1N343 N1N304 VDD VDD pch W=5.4U L=0.24U
M10 N1N343 N1N413 N1N345 VDD pch W=5.4U L=0.24U
M11 N1N345 N1N304 VSS VSS nch W=1.5U L=0.24U
M12 VSS N1N413 N1N345 VSS nch W=1.5U L=0.24U
M13 N1N413 DIN5 VDD VDD pch W=2.1U L=0.24U
M14 N1N413 DIN6 VDD VDD pch W=2.1U L=0.24U
M15 N1N413 DIN7 VDD VDD pch W=2.1U L=0.24U
M16 N1N413 DIN8 VDD VDD pch W=2.1U L=0.24U
M17 N1N413 DIN5 N1N362 VSS nch W=6.3U L=0.24U
M18 N1N362 DIN6 N1N364 VSS nch W=6.5U L=0.24U
M19 N1N364 DIN7 N1N366 VSS nch W=6.7U L=0.24U
M20 N1N366 DIN8 VSS VSS nch W=6.9U L=0.24U
M22 Q N1N345 VSS VSS nch W=3U L=0.24U
M21 Q N1N345 VDD VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nor2s1 Q DIN1 DIN2
M3 Q DIN1 VSS VSS nch W=0.7U L=0.24U
M1 N1N427 DIN1 VDD VDD pch W=3U L=0.24U
M2 Q DIN2 N1N427 VDD pch W=3U L=0.24U
M4 Q DIN2 VSS VSS nch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor Q DIN1 DIN2
M3 Q DIN1 VSS VSS nch W=0.7U L=0.24U
M1 N1N427 DIN1 VDD VDD pch W=3U L=0.24U
M2 Q DIN2 N1N427 VDD pch W=3U L=0.24U
M4 Q DIN2 VSS VSS nch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor2s2 Q DIN1 DIN2
M3 Q DIN1 VSS VSS nch W=1.5U L=0.24U
M1 N1N427 DIN1 VDD VDD pch W=6.34U L=0.24U
M2 Q DIN2 N1N427 VDD pch W=6.34U L=0.24U
M4 Q DIN2 VSS VSS nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor2s3 Q DIN1 DIN2
M3 Q DIN1 VSS VSS nch W=2.7U L=0.24U
M1 N1N427 DIN1 VDD VDD pch W=10.9U L=0.24U
M2 Q DIN2 N1N427 VDD pch W=10.9U L=0.24U
M4 Q DIN2 VSS VSS nch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor3s1 Q DIN1 DIN2 DIN3
M4 Q DIN1 VSS VSS nch W=0.74U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=4.38U L=0.24U
M2 N1N430 DIN2 N1N428 VDD pch W=4.38U L=0.24U
M3 Q DIN3 N1N430 VDD pch W=4.38U L=0.24U
M5 Q DIN2 VSS VSS nch W=0.74U L=0.24U
M6 Q DIN3 VSS VSS nch W=0.74U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor3s2 Q DIN1 DIN2 DIN3
M4 Q DIN1 VSS VSS nch W=1.7U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=9.4U L=0.24U
M2 N1N430 DIN2 N1N428 VDD pch W=9.4U L=0.24U
M3 Q DIN3 N1N430 VDD pch W=9.4U L=0.24U
M5 Q DIN2 VSS VSS nch W=1.7U L=0.24U
M6 Q DIN3 VSS VSS nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor3s3 Q DIN1 DIN2 DIN3
M4 Q DIN1 VSS VSS nch W=3.1U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=16U L=0.24U
M2 N1N430 DIN2 N1N428 VDD pch W=16U L=0.24U
M3 Q DIN3 N1N430 VDD pch W=16U L=0.24U
M5 Q DIN2 VSS VSS nch W=3.1U L=0.24U
M6 Q DIN3 VSS VSS nch W=3.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xor4s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 VSS VSS nch W=0.86U L=0.24U
M1 N1N452 DIN1 VDD VDD pch W=6.2U L=0.24U
M2 N1N450 DIN2 N1N452 VDD pch W=6U L=0.24U
M3 N1N448 DIN3 N1N450 VDD pch W=5.8U L=0.24U
M4 Q DIN4 N1N448 VDD pch W=5.5U L=0.24U
M6 Q DIN2 VSS VSS nch W=0.86U L=0.24U
M7 Q DIN3 VSS VSS nch W=0.86U L=0.24U
M8 Q DIN4 VSS VSS nch W=0.86U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xnr4s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 VSS VSS nch W=0.86U L=0.24U
M1 N1N452 DIN1 VDD VDD pch W=6.2U L=0.24U
M2 N1N450 DIN2 N1N452 VDD pch W=6U L=0.24U
M3 N1N448 DIN3 N1N450 VDD pch W=5.8U L=0.24U
M4 Q DIN4 N1N448 VDD pch W=5.5U L=0.24U
M6 Q DIN2 VSS VSS nch W=0.86U L=0.24U
M7 Q DIN3 VSS VSS nch W=0.86U L=0.24U
M8 Q DIN4 VSS VSS nch W=0.86U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nor4s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 VSS VSS nch W=0.86U L=0.24U
M1 N1N452 DIN1 VDD VDD pch W=6.2U L=0.24U
M2 N1N450 DIN2 N1N452 VDD pch W=6U L=0.24U
M3 N1N448 DIN3 N1N450 VDD pch W=5.8U L=0.24U
M4 Q DIN4 N1N448 VDD pch W=5.5U L=0.24U
M6 Q DIN2 VSS VSS nch W=0.86U L=0.24U
M7 Q DIN3 VSS VSS nch W=0.86U L=0.24U
M8 Q DIN4 VSS VSS nch W=0.86U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor4s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 VSS VSS nch W=1.7U L=0.24U
M1 N1N452 DIN1 VDD VDD pch W=12U L=0.24U
M2 N1N450 DIN2 N1N452 VDD pch W=11.8U L=0.24U
M3 N1N448 DIN3 N1N450 VDD pch W=11.4U L=0.24U
M4 Q DIN4 N1N448 VDD pch W=10.6U L=0.24U
M6 Q DIN2 VSS VSS nch W=1.7U L=0.24U
M7 Q DIN3 VSS VSS nch W=1.7U L=0.24U
M8 Q DIN4 VSS VSS nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor4s3 Q DIN1 DIN2 DIN3 DIN4
M3 N1N438 DIN1 VSS VSS nch W=1.8U L=0.24U
M1 N1N436 DIN1 VDD VDD pch W=5.2U L=0.24U
M2 N1N438 DIN2 N1N436 VDD pch W=4.4U L=0.24U
M4 N1N438 DIN2 VSS VSS nch W=1.8U L=0.24U
M5 N1N450 N1N438 VDD VDD pch W=4.2U L=0.24U
M6 VDD N1N457 N1N450 VDD pch W=3.8U L=0.24U
M7 N1N450 N1N438 N1N453 VSS nch W=4.4U L=0.24U
M8 N1N453 N1N457 VSS VSS nch W=4.4U L=0.24U
M9 N1N455 DIN3 VDD VDD pch W=5.2U L=0.24U
M10 N1N457 DIN4 N1N455 VDD pch W=4.4U L=0.24U
M11 N1N457 DIN3 VSS VSS nch W=1.8U L=0.24U
M12 N1N457 DIN4 VSS VSS nch W=1.8U L=0.24U
M14 Q N1N450 VSS VSS nch W=4.2U L=0.24U
M13 Q N1N450 VDD VDD pch W=8.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xor5s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 VSS VSS nch W=0.7U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=3.1U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=2.8U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=2.5U L=0.24U
M4 N1N444 DIN3 VSS VSS nch W=0.7U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=0.7U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=1.9U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=1.7U L=0.24U
M9 N1N494 DIN5 VSS VSS nch W=0.7U L=0.24U
M10 VSS DIN4 N1N494 VSS nch W=0.7U L=0.24U
M11 N1N474 N1N444 VDD VDD pch W=2U L=0.24U
M12 VDD N1N494 N1N474 VDD pch W=2U L=0.24U
M13 N1N474 N1N444 N1N480 VSS nch W=1.6U L=0.24U
M14 N1N480 N1N494 VSS VSS nch W=1.6U L=0.24U
M16 Q N1N474 VSS VSS nch W=1.1U L=0.24U
M15 Q N1N474 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT xnr5s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 VSS VSS nch W=0.7U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=3.1U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=2.8U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=2.5U L=0.24U
M4 N1N444 DIN3 VSS VSS nch W=0.7U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=0.7U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=1.9U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=1.7U L=0.24U
M9 N1N494 DIN5 VSS VSS nch W=0.7U L=0.24U
M10 VSS DIN4 N1N494 VSS nch W=0.7U L=0.24U
M11 N1N474 N1N444 VDD VDD pch W=2U L=0.24U
M12 VDD N1N494 N1N474 VDD pch W=2U L=0.24U
M13 N1N474 N1N444 N1N480 VSS nch W=1.6U L=0.24U
M14 N1N480 N1N494 VSS VSS nch W=1.6U L=0.24U
M16 Q N1N474 VSS VSS nch W=1.1U L=0.24U
M15 Q N1N474 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nor5s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 VSS VSS nch W=0.7U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=3.1U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=2.8U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=2.5U L=0.24U
M4 N1N444 DIN3 VSS VSS nch W=0.7U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=0.7U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=1.9U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=1.7U L=0.24U
M9 N1N494 DIN5 VSS VSS nch W=0.7U L=0.24U
M10 VSS DIN4 N1N494 VSS nch W=0.7U L=0.24U
M11 N1N474 N1N444 VDD VDD pch W=2U L=0.24U
M12 VDD N1N494 N1N474 VDD pch W=2U L=0.24U
M13 N1N474 N1N444 N1N480 VSS nch W=1.6U L=0.24U
M14 N1N480 N1N494 VSS VSS nch W=1.6U L=0.24U
M16 Q N1N474 VSS VSS nch W=1.1U L=0.24U
M15 Q N1N474 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor5s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 VSS VSS nch W=1.4U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=6.1U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=5.9U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=5.7U L=0.24U
M4 N1N444 DIN3 VSS VSS nch W=1.4U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=1.4U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=4U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=3.8U L=0.24U
M9 N1N494 DIN5 VSS VSS nch W=1.4U L=0.24U
M10 VSS DIN4 N1N494 VSS nch W=1.4U L=0.24U
M11 N1N474 N1N444 VDD VDD pch W=3.9U L=0.24U
M12 VDD N1N494 N1N474 VDD pch W=3.9U L=0.24U
M13 N1N474 N1N444 N1N480 VSS nch W=3.7U L=0.24U
M14 N1N480 N1N494 VSS VSS nch W=3.8U L=0.24U
M16 Q N1N474 VSS VSS nch W=2.1U L=0.24U
M15 Q N1N474 VDD VDD pch W=4.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor5s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 VSS VSS nch W=2.3U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=10.7U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=10.2U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=9.5U L=0.24U
M4 N1N444 DIN3 VSS VSS nch W=2.3U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=2.3U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=6.3U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=6.2U L=0.24U
M9 N1N494 DIN5 VSS VSS nch W=2.3U L=0.24U
M10 VSS DIN4 N1N494 VSS nch W=2.3U L=0.24U
M11 N1N474 N1N444 VDD VDD pch W=6.8U L=0.24U
M12 VDD N1N494 N1N474 VDD pch W=6.8U L=0.24U
M13 N1N474 N1N444 N1N480 VSS nch W=5.8U L=0.24U
M14 N1N480 N1N494 VSS VSS nch W=5.9U L=0.24U
M16 Q N1N474 VSS VSS nch W=4U L=0.24U
M15 Q N1N474 VDD VDD pch W=8.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xnr6s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M3 N1N421 DIN3 N1N425 VDD pch W=2.5U L=0.24U
M2 N1N425 DIN2 N1N426 VDD pch W=2.8U L=0.24U
M4 N1N421 DIN3 VSS VSS nch W=0.7U L=0.24U
M1 N1N426 DIN1 VDD VDD pch W=3.1U L=0.24U
M5 N1N421 DIN2 VSS VSS nch W=0.7U L=0.24U
M6 N1N421 DIN1 VSS VSS nch W=0.7U L=0.24U
M11 N1N428 DIN4 VDD VDD pch W=3.1U L=0.24U
M12 N1N423 DIN5 N1N428 VDD pch W=2.8U L=0.24U
M13 N1N434 DIN6 N1N423 VDD pch W=2.5U L=0.24U
M14 N1N434 DIN6 VSS VSS nch W=0.7U L=0.24U
M8 VDD N1N434 N1N453 VDD pch W=2U L=0.24U
M9 N1N453 N1N421 N1N451 VSS nch W=1.6U L=0.24U
M10 N1N451 N1N434 VSS VSS nch W=1.6U L=0.24U
M16 N1N434 DIN4 VSS VSS nch W=0.7U L=0.24U
M15 N1N434 DIN5 VSS VSS nch W=0.7U L=0.24U
M7 N1N453 N1N421 VDD VDD pch W=2U L=0.24U
M18 Q N1N453 VSS VSS nch W=1.1U L=0.24U
M17 Q N1N453 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT xor6s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M3 N1N421 DIN3 N1N425 VDD pch W=2.5U L=0.24U
M2 N1N425 DIN2 N1N426 VDD pch W=2.8U L=0.24U
M4 N1N421 DIN3 VSS VSS nch W=0.7U L=0.24U
M1 N1N426 DIN1 VDD VDD pch W=3.1U L=0.24U
M5 N1N421 DIN2 VSS VSS nch W=0.7U L=0.24U
M6 N1N421 DIN1 VSS VSS nch W=0.7U L=0.24U
M11 N1N428 DIN4 VDD VDD pch W=3.1U L=0.24U
M12 N1N423 DIN5 N1N428 VDD pch W=2.8U L=0.24U
M13 N1N434 DIN6 N1N423 VDD pch W=2.5U L=0.24U
M14 N1N434 DIN6 VSS VSS nch W=0.7U L=0.24U
M8 VDD N1N434 N1N453 VDD pch W=2U L=0.24U
M9 N1N453 N1N421 N1N451 VSS nch W=1.6U L=0.24U
M10 N1N451 N1N434 VSS VSS nch W=1.6U L=0.24U
M16 N1N434 DIN4 VSS VSS nch W=0.7U L=0.24U
M15 N1N434 DIN5 VSS VSS nch W=0.7U L=0.24U
M7 N1N453 N1N421 VDD VDD pch W=2U L=0.24U
M18 Q N1N453 VSS VSS nch W=1.1U L=0.24U
M17 Q N1N453 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT or6s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M3 N1N421 DIN3 N1N425 VDD pch W=2.5U L=0.24U
M2 N1N425 DIN2 N1N426 VDD pch W=2.8U L=0.24U
M4 N1N421 DIN3 VSS VSS nch W=0.7U L=0.24U
M1 N1N426 DIN1 VDD VDD pch W=3.1U L=0.24U
M5 N1N421 DIN2 VSS VSS nch W=0.7U L=0.24U
M6 N1N421 DIN1 VSS VSS nch W=0.7U L=0.24U
M11 N1N428 DIN4 VDD VDD pch W=3.1U L=0.24U
M12 N1N423 DIN5 N1N428 VDD pch W=2.8U L=0.24U
M13 N1N434 DIN6 N1N423 VDD pch W=2.5U L=0.24U
M14 N1N434 DIN6 VSS VSS nch W=0.7U L=0.24U
M8 VDD N1N434 N1N453 VDD pch W=2U L=0.24U
M9 N1N453 N1N421 N1N451 VSS nch W=1.6U L=0.24U
M10 N1N451 N1N434 VSS VSS nch W=1.6U L=0.24U
M16 N1N434 DIN4 VSS VSS nch W=0.7U L=0.24U
M15 N1N434 DIN5 VSS VSS nch W=0.7U L=0.24U
M7 N1N453 N1N421 VDD VDD pch W=2U L=0.24U
M18 Q N1N453 VSS VSS nch W=1.1U L=0.24U
M17 Q N1N453 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nor6s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M3 N1N421 DIN3 N1N425 VDD pch W=2.5U L=0.24U
M2 N1N425 DIN2 N1N426 VDD pch W=2.8U L=0.24U
M4 N1N421 DIN3 VSS VSS nch W=0.7U L=0.24U
M1 N1N426 DIN1 VDD VDD pch W=3.1U L=0.24U
M5 N1N421 DIN2 VSS VSS nch W=0.7U L=0.24U
M6 N1N421 DIN1 VSS VSS nch W=0.7U L=0.24U
M11 N1N428 DIN4 VDD VDD pch W=3.1U L=0.24U
M12 N1N423 DIN5 N1N428 VDD pch W=2.8U L=0.24U
M13 N1N434 DIN6 N1N423 VDD pch W=2.5U L=0.24U
M14 N1N434 DIN6 VSS VSS nch W=0.7U L=0.24U
M8 VDD N1N434 N1N453 VDD pch W=2U L=0.24U
M9 N1N453 N1N421 N1N451 VSS nch W=1.6U L=0.24U
M10 N1N451 N1N434 VSS VSS nch W=1.6U L=0.24U
M16 N1N434 DIN4 VSS VSS nch W=0.7U L=0.24U
M15 N1N434 DIN5 VSS VSS nch W=0.7U L=0.24U
M7 N1N453 N1N421 VDD VDD pch W=2U L=0.24U
M18 Q N1N453 VSS VSS nch W=1.1U L=0.24U
M17 Q N1N453 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor6s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N444 DIN3 VSS VSS nch W=1.4U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=6.1U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=5.9U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=5.7U L=0.24U
M11 N1N460 DIN4 VDD VDD pch W=6.1U L=0.24U
M5 N1N444 DIN2 VSS VSS nch W=1.4U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=1.4U L=0.24U
M12 N1N462 DIN5 N1N460 VDD pch W=5.9U L=0.24U
M13 N1N464 DIN6 N1N462 VDD pch W=5.7U L=0.24U
M14 N1N464 DIN6 VSS VSS nch W=1.4U L=0.24U
M15 N1N464 DIN5 VSS VSS nch W=1.4U L=0.24U
M16 N1N464 DIN4 VSS VSS nch W=1.4U L=0.24U
M7 N1N480 N1N444 VDD VDD pch W=3.9U L=0.24U
M8 VDD N1N464 N1N480 VDD pch W=3.9U L=0.24U
M9 N1N480 N1N444 N1N483 VSS nch W=3.7U L=0.24U
M10 N1N483 N1N464 VSS VSS nch W=3.8U L=0.24U
M18 Q N1N480 VSS VSS nch W=2.1U L=0.24U
M17 Q N1N480 VDD VDD pch W=4.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT nor6s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N506 DIN3 VSS VSS nch W=2.3U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=10.7U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=10.2U L=0.24U
M3 N1N506 DIN3 N1N442 VDD pch W=9.5U L=0.24U
M11 N1N460 DIN4 VDD VDD pch W=10.7U L=0.24U
M5 N1N506 DIN2 VSS VSS nch W=2.3U L=0.24U
M6 N1N506 DIN1 VSS VSS nch W=2.3U L=0.24U
M12 N1N462 DIN5 N1N460 VDD pch W=10.2U L=0.24U
M13 N1N464 DIN6 N1N462 VDD pch W=9.5U L=0.24U
M14 N1N464 DIN6 VSS VSS nch W=2.3U L=0.24U
M15 N1N464 DIN5 VSS VSS nch W=2.3U L=0.24U
M16 N1N464 DIN4 VSS VSS nch W=2.3U L=0.24U
M7 N1N480 N1N506 VDD VDD pch W=6.8U L=0.24U
M8 VDD N1N464 N1N480 VDD pch W=6.8U L=0.24U
M9 N1N480 N1N506 N1N483 VSS nch W=5.8U L=0.24U
M10 N1N483 N1N464 VSS VSS nch W=5.9U L=0.24U
M18 Q N1N480 VSS VSS nch W=4U L=0.24U
M17 Q N1N480 VDD VDD pch W=8.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or7s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M4 N1N446 DIN1 VSS VSS nch W=2.34U L=0.24U
M1 N1N441 DIN1 VDD VDD pch W=9U L=0.24U
M2 N1N443 DIN2 N1N441 VDD pch W=8.8U L=0.24U
M3 N1N446 DIN3 N1N443 VDD pch W=8.6U L=0.24U
M5 N1N446 DIN2 VSS VSS nch W=2.34U L=0.24U
M6 N1N446 DIN3 VSS VSS nch W=2.34U L=0.24U
M7 N1N465 N1N446 VDD VDD pch W=5.4U L=0.24U
M8 VDD N1N471 N1N465 VDD pch W=5.4U L=0.24U
M9 N1N465 N1N446 N1N473 VSS nch W=5U L=0.24U
M10 VSS N1N471 N1N473 VSS nch W=5U L=0.24U
M11 N1N478 DIN4 VDD VDD pch W=11.7U L=0.24U
M12 N1N480 DIN5 N1N478 VDD pch W=11.5U L=0.24U
M13 N1N491 DIN6 N1N480 VDD pch W=11.3U L=0.24U
M16 N1N471 DIN6 VSS VSS nch W=2.34U L=0.24U
M17 N1N471 DIN5 VSS VSS nch W=2.34U L=0.24U
M18 N1N471 DIN4 VSS VSS nch W=2.34U L=0.24U
M15 N1N471 DIN7 VSS VSS nch W=2.34U L=0.24U
M14 N1N471 DIN7 N1N491 VDD pch W=11.1U L=0.24U
M19 Q N1N465 VDD VDD pch W=7U L=0.24U
M20 Q N1N465 VSS VSS nch W=3.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT xor7s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M4 N1N446 DIN1 VSS VSS nch W=2.34U L=0.24U
M1 N1N441 DIN1 VDD VDD pch W=9U L=0.24U
M2 N1N443 DIN2 N1N441 VDD pch W=8.8U L=0.24U
M3 N1N446 DIN3 N1N443 VDD pch W=8.6U L=0.24U
M5 N1N446 DIN2 VSS VSS nch W=2.34U L=0.24U
M6 N1N446 DIN3 VSS VSS nch W=2.34U L=0.24U
M7 N1N465 N1N446 VDD VDD pch W=5.4U L=0.24U
M8 VDD N1N471 N1N465 VDD pch W=5.4U L=0.24U
M9 N1N465 N1N446 N1N473 VSS nch W=5U L=0.24U
M10 VSS N1N471 N1N473 VSS nch W=5U L=0.24U
M11 N1N478 DIN4 VDD VDD pch W=11.7U L=0.24U
M12 N1N480 DIN5 N1N478 VDD pch W=11.5U L=0.24U
M13 N1N491 DIN6 N1N480 VDD pch W=11.3U L=0.24U
M16 N1N471 DIN6 VSS VSS nch W=2.34U L=0.24U
M17 N1N471 DIN5 VSS VSS nch W=2.34U L=0.24U
M18 N1N471 DIN4 VSS VSS nch W=2.34U L=0.24U
M15 N1N471 DIN7 VSS VSS nch W=2.34U L=0.24U
M14 N1N471 DIN7 N1N491 VDD pch W=11.1U L=0.24U
M19 Q N1N465 VDD VDD pch W=7U L=0.24U
M20 Q N1N465 VSS VSS nch W=3.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT xnr7s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M4 N1N446 DIN1 VSS VSS nch W=2.34U L=0.24U
M1 N1N441 DIN1 VDD VDD pch W=9U L=0.24U
M2 N1N443 DIN2 N1N441 VDD pch W=8.8U L=0.24U
M3 N1N446 DIN3 N1N443 VDD pch W=8.6U L=0.24U
M5 N1N446 DIN2 VSS VSS nch W=2.34U L=0.24U
M6 N1N446 DIN3 VSS VSS nch W=2.34U L=0.24U
M7 N1N465 N1N446 VDD VDD pch W=5.4U L=0.24U
M8 VDD N1N471 N1N465 VDD pch W=5.4U L=0.24U
M9 N1N465 N1N446 N1N473 VSS nch W=5U L=0.24U
M10 VSS N1N471 N1N473 VSS nch W=5U L=0.24U
M11 N1N478 DIN4 VDD VDD pch W=11.7U L=0.24U
M12 N1N480 DIN5 N1N478 VDD pch W=11.5U L=0.24U
M13 N1N491 DIN6 N1N480 VDD pch W=11.3U L=0.24U
M16 N1N471 DIN6 VSS VSS nch W=2.34U L=0.24U
M17 N1N471 DIN5 VSS VSS nch W=2.34U L=0.24U
M18 N1N471 DIN4 VSS VSS nch W=2.34U L=0.24U
M15 N1N471 DIN7 VSS VSS nch W=2.34U L=0.24U
M14 N1N471 DIN7 N1N491 VDD pch W=11.1U L=0.24U
M19 Q N1N465 VDD VDD pch W=7U L=0.24U
M20 Q N1N465 VSS VSS nch W=3.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
.SUBCKT nor7s3 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M4 N1N446 DIN1 VSS VSS nch W=2.34U L=0.24U
M1 N1N441 DIN1 VDD VDD pch W=9U L=0.24U
M2 N1N443 DIN2 N1N441 VDD pch W=8.8U L=0.24U
M3 N1N446 DIN3 N1N443 VDD pch W=8.6U L=0.24U
M5 N1N446 DIN2 VSS VSS nch W=2.34U L=0.24U
M6 N1N446 DIN3 VSS VSS nch W=2.34U L=0.24U
M7 N1N465 N1N446 VDD VDD pch W=5.4U L=0.24U
M8 VDD N1N471 N1N465 VDD pch W=5.4U L=0.24U
M9 N1N465 N1N446 N1N473 VSS nch W=5U L=0.24U
M10 VSS N1N471 N1N473 VSS nch W=5U L=0.24U
M11 N1N478 DIN4 VDD VDD pch W=11.7U L=0.24U
M12 N1N480 DIN5 N1N478 VDD pch W=11.5U L=0.24U
M13 N1N491 DIN6 N1N480 VDD pch W=11.3U L=0.24U
M16 N1N471 DIN6 VSS VSS nch W=2.34U L=0.24U
M17 N1N471 DIN5 VSS VSS nch W=2.34U L=0.24U
M18 N1N471 DIN4 VSS VSS nch W=2.34U L=0.24U
M15 N1N471 DIN7 VSS VSS nch W=2.34U L=0.24U
M14 N1N471 DIN7 N1N491 VDD pch W=11.1U L=0.24U
M19 Q N1N465 VDD VDD pch W=7U L=0.24U
M20 Q N1N465 VSS VSS nch W=3.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT npd1s1 OUTD GIN
M1 OUTD GIN VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT npd1s2 OUTD GIN
M1 OUTD GIN VSS VSS nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT npt1s1 DIN OUTD OUTS
M1 OUTD DIN OUTS VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT npt1s2 DIN OUTD OUTS
M1 OUTD DIN OUTS VSS nch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT npt1s3 DIN OUTD OUTS
M1 OUTD DIN OUTS VSS nch W=8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT npt1s4 DIN OUTD OUTS
M1 OUTD DIN OUTS VSS nch W=16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT npt1s5 DIN OUTD OUTS
M1 OUTD DIN OUTS VSS nch W=32U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT npt1s6 DIN OUTS OUTD
M1 OUTD DIN OUTS VSS nch W=65U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oaaoi1123s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 Q DIN7 VSS VSS nch W=0.6U L=0.24U
M7 Q DIN7 N1N349 VDD pch W=6.9U L=0.24U
M4 N1N349 DIN6 N1N360 VDD pch W=6.9U L=0.24U
M5 N1N360 DIN4 N1N283 VDD pch W=6.9U L=0.24U
M6 N1N349 DIN5 N1N283 VDD pch W=6.9U L=0.24U
M3 VDD DIN3 N1N360 VDD pch W=6.9U L=0.24U
M1 N1N360 DIN2 VDD VDD pch W=6.9U L=0.24U
M2 N1N360 DIN1 VDD VDD pch W=6.9U L=0.24U
M9 Q DIN6 N1N315 VSS nch W=1U L=0.24U
M10 N1N289 DIN3 Q VSS nch W=1.3U L=0.24U
M12 N1N315 DIN5 VSS VSS nch W=1U L=0.24U
M11 N1N315 DIN4 VSS VSS nch W=1U L=0.24U
M13 N1N289 DIN2 N1N291 VSS nch W=1.3U L=0.24U
M14 N1N291 DIN1 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oaaoi1123s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 N1N302 DIN7 VSS VSS nch W=0.6U L=0.24U
M7 N1N302 DIN7 N1N349 VDD pch W=6.9U L=0.24U
M4 N1N349 DIN6 N1N360 VDD pch W=6.9U L=0.24U
M5 N1N360 DIN4 N1N283 VDD pch W=6.9U L=0.24U
M6 N1N349 DIN5 N1N283 VDD pch W=6.9U L=0.24U
M3 VDD DIN3 N1N360 VDD pch W=6.9U L=0.24U
M1 N1N360 DIN2 VDD VDD pch W=6.9U L=0.24U
M2 N1N360 DIN1 VDD VDD pch W=6.9U L=0.24U
M9 N1N302 DIN6 N1N315 VSS nch W=1U L=0.24U
M10 N1N289 DIN3 N1N302 VSS nch W=1.3U L=0.24U
M12 N1N315 DIN5 VSS VSS nch W=1U L=0.24U
M11 N1N315 DIN4 VSS VSS nch W=1U L=0.24U
M13 N1N289 DIN2 N1N291 VSS nch W=1.3U L=0.24U
M14 N1N291 DIN1 VSS VSS nch W=1.3U L=0.24U
M15 N1N371 N1N302 VDD VDD pch W=3.7U L=0.24U
M16 N1N371 N1N302 VSS VSS nch W=1.6U L=0.24U
M18 Q N1N371 VSS VSS nch W=4.1U L=0.24U
M17 Q N1N371 VDD VDD pch W=7.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oaaoi1123s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 N1N302 DIN7 VSS VSS nch W=0.6U L=0.24U
M7 N1N302 DIN7 N1N349 VDD pch W=6.9U L=0.24U
M4 N1N349 DIN6 N1N360 VDD pch W=6.9U L=0.24U
M5 N1N360 DIN4 N1N283 VDD pch W=6.9U L=0.24U
M6 N1N349 DIN5 N1N283 VDD pch W=6.9U L=0.24U
M3 VDD DIN3 N1N360 VDD pch W=6.9U L=0.24U
M1 N1N360 DIN2 VDD VDD pch W=6.9U L=0.24U
M2 N1N360 DIN1 VDD VDD pch W=6.9U L=0.24U
M9 N1N302 DIN6 N1N315 VSS nch W=1U L=0.24U
M10 N1N289 DIN3 N1N302 VSS nch W=1.3U L=0.24U
M12 N1N315 DIN5 VSS VSS nch W=1U L=0.24U
M11 N1N315 DIN4 VSS VSS nch W=1U L=0.24U
M13 N1N289 DIN2 N1N291 VSS nch W=1.3U L=0.24U
M14 N1N291 DIN1 VSS VSS nch W=1.3U L=0.24U
M15 N1N371 N1N302 VDD VDD pch W=5.2U L=0.24U
M16 N1N371 N1N302 VSS VSS nch W=2.2U L=0.24U
M18 Q N1N371 VSS VSS nch W=5.7U L=0.24U
M17 Q N1N371 VDD VDD pch W=10.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai1112s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N284 VSS nch W=1.4U L=0.24U
M1 Q DIN1 VDD VDD pch W=0.7U L=0.24U
M2 Q DIN2 VDD VDD pch W=0.7U L=0.24U
M3 Q DIN3 VDD VDD pch W=0.7U L=0.24U
M4 VDD DIN4 N1N302 VDD pch W=1.4U L=0.24U
M5 N1N302 DIN5 Q VDD pch W=1.4U L=0.24U
M7 N1N284 DIN2 N1N286 VSS nch W=1.4U L=0.24U
M8 N1N286 DIN3 N1N292 VSS nch W=1.4U L=0.24U
M9 N1N292 DIN4 VSS VSS nch W=1.4U L=0.24U
M10 VSS DIN5 N1N292 VSS nch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai1112s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N284 VSS nch W=2U L=0.24U
M1 Q DIN1 VDD VDD pch W=1U L=0.24U
M2 Q DIN2 VDD VDD pch W=1U L=0.24U
M3 Q DIN3 VDD VDD pch W=1U L=0.24U
M4 VDD DIN4 N1N302 VDD pch W=2U L=0.24U
M5 N1N302 DIN5 Q VDD pch W=2U L=0.24U
M7 N1N284 DIN2 N1N286 VSS nch W=2U L=0.24U
M8 N1N286 DIN3 N1N292 VSS nch W=2U L=0.24U
M9 N1N292 DIN4 VSS VSS nch W=2U L=0.24U
M10 VSS DIN5 N1N292 VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai1112s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N278 DIN1 N1N284 VSS nch W=1.8U L=0.24U
M1 N1N278 DIN1 VDD VDD pch W=0.9U L=0.24U
M2 N1N278 DIN2 VDD VDD pch W=0.9U L=0.24U
M3 N1N278 DIN3 VDD VDD pch W=0.9U L=0.24U
M4 VDD DIN4 N1N302 VDD pch W=1.8U L=0.24U
M5 N1N302 DIN5 N1N278 VDD pch W=1.8U L=0.24U
M7 N1N284 DIN2 N1N286 VSS nch W=1.8U L=0.24U
M8 N1N286 DIN3 N1N292 VSS nch W=1.9U L=0.24U
M9 N1N292 DIN4 VSS VSS nch W=1.9U L=0.24U
M10 VSS DIN5 N1N292 VSS nch W=1.9U L=0.24U
M11 N1N326 N1N278 VDD VDD pch W=3.4U L=0.24U
M12 N1N326 N1N278 VSS VSS nch W=1.8U L=0.24U
M14 Q N1N326 VSS VSS nch W=3.1U L=0.24U
M13 Q N1N326 VDD VDD pch W=5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai13s1 Q DIN1 DIN2 DIN3 DIN4
M1 N1N330 DIN2 VDD VDD pch W=1.8U L=0.24U
M6 N1N339 DIN2 VSS VSS nch W=0.7U L=0.24U
M2 N1N332 DIN3 N1N330 VDD pch W=1.8U L=0.24U
M3 Q DIN4 N1N332 VDD pch W=1.8U L=0.24U
M4 VDD DIN1 Q VDD pch W=0.66U L=0.24U
M7 N1N339 DIN3 VSS VSS nch W=0.7U L=0.24U
M8 VSS DIN4 N1N339 VSS nch W=0.7U L=0.24U
M5 N1N339 DIN1 Q VSS nch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai13s2 Q DIN1 DIN2 DIN3 DIN4
M1 N1N330 DIN2 VDD VDD pch W=2.16U L=0.24U
M6 N1N339 DIN2 VSS VSS nch W=0.84U L=0.24U
M2 N1N332 DIN3 N1N330 VDD pch W=2.16U L=0.24U
M3 Q DIN4 N1N332 VDD pch W=2.16U L=0.24U
M4 VDD DIN1 Q VDD pch W=0.8U L=0.24U
M7 N1N339 DIN3 VSS VSS nch W=0.84U L=0.24U
M8 VSS DIN4 N1N339 VSS nch W=0.84U L=0.24U
M5 N1N339 DIN1 Q VSS nch W=0.84U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai13s3 Q DIN1 DIN2 DIN3 DIN4
M1 N1N330 DIN2 VDD VDD pch W=1.8U L=0.24U
M6 N1N339 DIN2 VSS VSS nch W=0.9U L=0.24U
M2 N1N332 DIN3 N1N330 VDD pch W=1.8U L=0.24U
M3 N1N334 DIN4 N1N332 VDD pch W=1.8U L=0.24U
M4 VDD DIN1 N1N334 VDD pch W=0.66U L=0.24U
M7 N1N339 DIN3 VSS VSS nch W=0.9U L=0.24U
M8 VSS DIN4 N1N339 VSS nch W=0.9U L=0.24U
M5 N1N339 DIN1 N1N334 VSS nch W=0.9U L=0.24U
M10 N1N383 N1N334 VSS VSS nch W=1.2U L=0.24U
M12 Q N1N383 VSS VSS nch W=2U L=0.24U
M9 N1N383 N1N334 VDD VDD pch W=2.3U L=0.24U
M11 Q N1N383 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai211s1 Q DIN1 DIN2 DIN3 DIN4
M6 N1N469 DIN3 N1N444 VSS nch W=0.8U L=0.24U
M1 N1N435 DIN1 VDD VDD pch W=1.8U L=0.24U
M2 Q DIN2 N1N435 VDD pch W=1.8U L=0.24U
M3 Q DIN3 VDD VDD pch W=0.7U L=0.24U
M4 VDD DIN4 Q VDD pch W=0.7U L=0.24U
M7 N1N444 DIN1 VSS VSS nch W=0.8U L=0.24U
M5 N1N469 DIN4 Q VSS nch W=0.7U L=0.24U
M8 VSS DIN2 N1N444 VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai211s2 Q DIN1 DIN2 DIN3 DIN4
M6 N1N469 DIN3 N1N444 VSS nch W=1.2U L=0.24U
M1 N1N435 DIN1 VDD VDD pch W=2.9U L=0.24U
M2 Q DIN2 N1N435 VDD pch W=2.8U L=0.24U
M3 Q DIN3 VDD VDD pch W=1.1U L=0.24U
M4 VDD DIN4 Q VDD pch W=1.1U L=0.24U
M7 N1N444 DIN1 VSS VSS nch W=1.3U L=0.24U
M5 N1N469 DIN4 Q VSS nch W=1.1U L=0.24U
M8 VSS DIN2 N1N444 VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai211s3 Q DIN1 DIN2 DIN3 DIN4
M6 N1N326 DIN3 N1N327 VSS nch W=0.9U L=0.24U
M1 N1N332 DIN1 VDD VDD pch W=2U L=0.24U
M2 N1N329 DIN2 N1N332 VDD pch W=2U L=0.24U
M3 N1N329 DIN3 VDD VDD pch W=0.8U L=0.24U
M4 VDD DIN4 N1N329 VDD pch W=0.8U L=0.24U
M7 N1N327 DIN1 VSS VSS nch W=0.9U L=0.24U
M5 N1N326 DIN4 N1N329 VSS nch W=0.8U L=0.24U
M8 VSS DIN2 N1N327 VSS nch W=0.9U L=0.24U
M10 N1N374 N1N329 VSS VSS nch W=1.2U L=0.24U
M9 N1N374 N1N329 VDD VDD pch W=2U L=0.24U
M11 Q N1N374 VDD VDD pch W=4.3U L=0.24U
M12 Q N1N374 VSS VSS nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai21s1 Q DIN1 DIN2 DIN3
M5 N1N261 DIN2 VSS VSS nch W=0.6U L=0.24U
M1 Q DIN3 VDD VDD pch W=0.7U L=0.24U
M2 VDD DIN1 N1N257 VDD pch W=1.7U L=0.24U
M3 N1N257 DIN2 Q VDD pch W=1.7U L=0.24U
M4 Q DIN3 N1N261 VSS nch W=0.6U L=0.24U
M6 VSS DIN1 N1N261 VSS nch W=0.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai21s2 Q DIN1 DIN2 DIN3
M5 N1N284 DIN2 VSS VSS nch W=1U L=0.24U
M1 Q DIN3 VDD VDD pch W=1.2U L=0.24U
M2 VDD DIN1 N1N257 VDD pch W=2.8U L=0.24U
M3 N1N257 DIN2 Q VDD pch W=2.7U L=0.24U
M4 Q DIN3 N1N284 VSS nch W=1U L=0.24U
M6 VSS DIN1 N1N284 VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai21s3 Q DIN1 DIN2 DIN3
M5 N1N284 DIN2 VSS VSS nch W=2U L=0.24U
M1 Q DIN3 VDD VDD pch W=2.1U L=0.24U
M2 VDD DIN1 N1N257 VDD pch W=5.6U L=0.24U
M3 N1N257 DIN2 Q VDD pch W=5.4U L=0.24U
M4 Q DIN3 N1N284 VSS nch W=2U L=0.24U
M6 VSS DIN1 N1N284 VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai221s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M7 N1N283 DIN3 N1N292 VSS nch W=0.8U L=0.24U
M1 N1N263 DIN1 VDD VDD pch W=1.8U L=0.24U
M2 Q DIN2 N1N263 VDD pch W=1.8U L=0.24U
M3 VDD DIN3 N1N290 VDD pch W=1.8U L=0.24U
M5 VDD DIN5 Q VDD pch W=0.8U L=0.24U
M4 N1N290 DIN4 Q VDD pch W=1.8U L=0.24U
M9 N1N292 DIN1 VSS VSS nch W=0.8U L=0.24U
M10 VSS DIN2 N1N292 VSS nch W=0.8U L=0.24U
M8 N1N292 DIN4 N1N283 VSS nch W=0.8U L=0.24U
M6 N1N283 DIN5 Q VSS nch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai221s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M7 N1N283 DIN3 N1N292 VSS nch W=1.2U L=0.24U
M1 N1N263 DIN1 VDD VDD pch W=2.9U L=0.24U
M2 Q DIN2 N1N263 VDD pch W=2.8U L=0.24U
M3 VDD DIN3 N1N290 VDD pch W=2.9U L=0.24U
M5 VDD DIN5 Q VDD pch W=1.1U L=0.24U
M4 N1N290 DIN4 Q VDD pch W=2.8U L=0.24U
M9 N1N292 DIN1 VSS VSS nch W=1.3U L=0.24U
M10 VSS DIN2 N1N292 VSS nch W=1.3U L=0.24U
M8 N1N292 DIN4 N1N283 VSS nch W=1.2U L=0.24U
M6 N1N283 DIN5 Q VSS nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai221s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M7 N1N283 DIN3 N1N292 VSS nch W=0.9U L=0.24U
M1 N1N263 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N265 DIN2 N1N263 VDD pch W=2U L=0.24U
M3 VDD DIN3 N1N290 VDD pch W=2.1U L=0.24U
M5 VDD DIN5 N1N265 VDD pch W=0.8U L=0.24U
M4 N1N290 DIN4 N1N265 VDD pch W=2U L=0.24U
M9 N1N292 DIN1 VSS VSS nch W=1U L=0.24U
M10 VSS DIN2 N1N292 VSS nch W=1U L=0.24U
M8 N1N292 DIN4 N1N283 VSS nch W=0.9U L=0.24U
M6 N1N283 DIN5 N1N265 VSS nch W=0.8U L=0.24U
M12 N1N351 N1N265 VSS VSS nch W=1.3U L=0.24U
M11 N1N351 N1N265 VDD VDD pch W=2.2U L=0.24U
M13 Q N1N351 VDD VDD pch W=4.5U L=0.24U
M14 Q N1N351 VSS VSS nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai2222s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8
M3 N1N271 DIN2 N1N273 VSS nch W=0.7U L=0.24U
M6 N1N271 DIN1 N1N276 VDD pch W=1U L=0.24U
M2 N1N271 DIN3 N1N269 VDD pch W=1U L=0.24U
M4 N1N273 DIN3 VSS VSS nch W=0.7U L=0.24U
M1 N1N269 DIN4 VDD VDD pch W=1U L=0.24U
M5 N1N276 DIN2 VDD VDD pch W=1U L=0.24U
M7 N1N271 DIN1 N1N273 VSS nch W=0.7U L=0.24U
M8 N1N273 DIN4 VSS VSS nch W=0.7U L=0.24U
M11 N1N315 DIN6 N1N319 VSS nch W=0.7U L=0.24U
M9 N1N354 DIN8 VDD VDD pch W=1U L=0.24U
M10 N1N315 DIN7 N1N354 VDD pch W=1U L=0.24U
M12 N1N319 DIN7 VSS VSS nch W=0.7U L=0.24U
M16 N1N319 DIN8 VSS VSS nch W=0.7U L=0.24U
M15 N1N315 DIN5 N1N319 VSS nch W=0.7U L=0.24U
M13 N1N325 DIN6 VDD VDD pch W=1U L=0.24U
M14 N1N315 DIN5 N1N325 VDD pch W=1U L=0.24U
M19 N1N328 N1N271 VSS VSS nch W=0.6U L=0.24U
M18 N1N328 N1N271 N1N357 VDD pch W=1.5U L=0.24U
M17 VDD N1N315 N1N357 VDD pch W=1.5U L=0.24U
M20 N1N328 N1N315 VSS VSS nch W=0.6U L=0.24U
M22 Q N1N328 VSS VSS nch W=1U L=0.24U
M21 Q N1N328 VDD VDD pch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai2222s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8
M3 N1N271 DIN2 N1N273 VSS nch W=0.7U L=0.24U
M6 N1N271 DIN1 N1N276 VDD pch W=1U L=0.24U
M2 N1N271 DIN3 N1N269 VDD pch W=1U L=0.24U
M4 N1N273 DIN3 VSS VSS nch W=0.7U L=0.24U
M1 N1N269 DIN4 VDD VDD pch W=1U L=0.24U
M5 N1N276 DIN2 VDD VDD pch W=1U L=0.24U
M7 N1N271 DIN1 N1N273 VSS nch W=0.7U L=0.24U
M8 N1N273 DIN4 VSS VSS nch W=0.7U L=0.24U
M11 N1N315 DIN6 N1N319 VSS nch W=0.7U L=0.24U
M9 N1N354 DIN8 VDD VDD pch W=1U L=0.24U
M10 N1N315 DIN7 N1N354 VDD pch W=1U L=0.24U
M12 N1N319 DIN7 VSS VSS nch W=0.7U L=0.24U
M16 N1N319 DIN8 VSS VSS nch W=0.7U L=0.24U
M15 N1N315 DIN5 N1N319 VSS nch W=0.7U L=0.24U
M13 N1N325 DIN6 VDD VDD pch W=1U L=0.24U
M14 N1N315 DIN5 N1N325 VDD pch W=1U L=0.24U
M19 N1N328 N1N271 VSS VSS nch W=0.9U L=0.24U
M18 N1N328 N1N271 N1N357 VDD pch W=2.2U L=0.24U
M17 VDD N1N315 N1N357 VDD pch W=2.2U L=0.24U
M20 N1N328 N1N315 VSS VSS nch W=0.9U L=0.24U
M22 Q N1N328 VSS VSS nch W=1.4U L=0.24U
M21 Q N1N328 VDD VDD pch W=3.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai2222s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8
M3 N1N271 DIN2 N1N273 VSS nch W=1.4U L=0.24U
M6 N1N271 DIN1 N1N276 VDD pch W=2U L=0.24U
M2 N1N271 DIN3 N1N269 VDD pch W=2U L=0.24U
M4 N1N273 DIN3 VSS VSS nch W=1.4U L=0.24U
M1 N1N269 DIN4 VDD VDD pch W=2U L=0.24U
M5 N1N276 DIN2 VDD VDD pch W=2U L=0.24U
M7 N1N271 DIN1 N1N273 VSS nch W=1.4U L=0.24U
M8 N1N273 DIN4 VSS VSS nch W=1.4U L=0.24U
M11 N1N315 DIN6 N1N319 VSS nch W=1.4U L=0.24U
M9 N1N354 DIN8 VDD VDD pch W=2U L=0.24U
M10 N1N315 DIN7 N1N354 VDD pch W=2U L=0.24U
M12 N1N319 DIN7 VSS VSS nch W=1.4U L=0.24U
M16 N1N319 DIN8 VSS VSS nch W=1.4U L=0.24U
M15 N1N315 DIN5 N1N319 VSS nch W=1.4U L=0.24U
M13 N1N325 DIN6 VDD VDD pch W=2U L=0.24U
M14 N1N315 DIN5 N1N325 VDD pch W=2U L=0.24U
M19 N1N328 N1N271 VSS VSS nch W=1.5U L=0.24U
M18 N1N328 N1N271 N1N357 VDD pch W=3.4U L=0.24U
M17 VDD N1N315 N1N357 VDD pch W=3.4U L=0.24U
M20 N1N328 N1N315 VSS VSS nch W=1.5U L=0.24U
M22 Q N1N328 VSS VSS nch W=2.1U L=0.24U
M21 Q N1N328 VDD VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai222s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN5 N1N334 VSS nch W=0.9U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=1.9U L=0.24U
M4 Q DIN2 N1N323 VDD pch W=1.9U L=0.24U
M2 VDD DIN3 N1N325 VDD pch W=1.9U L=0.24U
M5 N1N325 DIN4 Q VDD pch W=1.9U L=0.24U
M3 VDD DIN5 N1N327 VDD pch W=1.9U L=0.24U
M6 N1N327 DIN6 Q VDD pch W=1.9U L=0.24U
M9 N1N334 DIN3 N1N338 VSS nch W=0.9U L=0.24U
M11 N1N338 DIN1 VSS VSS nch W=0.9U L=0.24U
M12 VSS DIN2 N1N338 VSS nch W=0.9U L=0.24U
M10 N1N338 DIN4 N1N334 VSS nch W=0.9U L=0.24U
M8 N1N334 DIN6 Q VSS nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai222s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N329 DIN5 N1N334 VSS nch W=0.9U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=2U L=0.24U
M4 N1N329 DIN2 N1N323 VDD pch W=1.9U L=0.24U
M2 VDD DIN3 N1N325 VDD pch W=2U L=0.24U
M5 N1N325 DIN4 N1N329 VDD pch W=1.9U L=0.24U
M3 VDD DIN5 N1N327 VDD pch W=2U L=0.24U
M6 N1N327 DIN6 N1N329 VDD pch W=1.9U L=0.24U
M9 N1N334 DIN3 N1N338 VSS nch W=0.9U L=0.24U
M11 N1N338 DIN1 VSS VSS nch W=1U L=0.24U
M12 VSS DIN2 N1N338 VSS nch W=1U L=0.24U
M10 N1N338 DIN4 N1N334 VSS nch W=0.9U L=0.24U
M8 N1N334 DIN6 N1N329 VSS nch W=0.9U L=0.24U
M14 N1N370 N1N329 VSS VSS nch W=0.6U L=0.24U
M13 N1N370 N1N329 VDD VDD pch W=1.3U L=0.24U
M15 Q N1N370 VDD VDD pch W=2.4U L=0.24U
M16 Q N1N370 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai222s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N329 DIN5 N1N334 VSS nch W=0.9U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=2.04U L=0.24U
M4 N1N329 DIN2 N1N323 VDD pch W=1.9U L=0.24U
M2 VDD DIN3 N1N325 VDD pch W=2.04U L=0.24U
M5 N1N325 DIN4 N1N329 VDD pch W=1.9U L=0.24U
M3 VDD DIN5 N1N327 VDD pch W=2.04U L=0.24U
M6 N1N327 DIN6 N1N329 VDD pch W=1.9U L=0.24U
M9 N1N334 DIN3 N1N338 VSS nch W=1U L=0.24U
M11 N1N338 DIN1 VSS VSS nch W=1.1U L=0.24U
M12 VSS DIN2 N1N338 VSS nch W=1.1U L=0.24U
M10 N1N338 DIN4 N1N334 VSS nch W=1U L=0.24U
M8 N1N334 DIN6 N1N329 VSS nch W=0.9U L=0.24U
M14 N1N372 N1N329 VSS VSS nch W=1U L=0.24U
M13 N1N372 N1N329 VDD VDD pch W=2.2U L=0.24U
M16 Q N1N372 VSS VSS nch W=2.1U L=0.24U
M15 Q N1N372 VDD VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai22s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N278 VSS nch W=0.64U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=1.7U L=0.24U
M2 Q DIN2 N1N258 VDD pch W=1.7U L=0.24U
M4 N1N260 DIN4 Q VDD pch W=1.7U L=0.24U
M3 VDD DIN3 N1N260 VDD pch W=1.7U L=0.24U
M6 N1N278 DIN3 VSS VSS nch W=0.64U L=0.24U
M8 VSS DIN4 N1N278 VSS nch W=0.64U L=0.24U
M7 N1N278 DIN2 Q VSS nch W=0.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai22s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N278 VSS nch W=1.02U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=2.6U L=0.24U
M2 Q DIN2 N1N258 VDD pch W=2.6U L=0.24U
M4 N1N260 DIN4 Q VDD pch W=2.6U L=0.24U
M3 VDD DIN3 N1N260 VDD pch W=2.6U L=0.24U
M6 N1N278 DIN3 VSS VSS nch W=1.02U L=0.24U
M8 VSS DIN4 N1N278 VSS nch W=1.02U L=0.24U
M7 N1N278 DIN2 Q VSS nch W=1.02U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai22s3 Q DIN1 DIN2 DIN3 DIN4
M5 N1N268 DIN1 N1N278 VSS nch W=0.8U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=1.8U L=0.24U
M2 N1N268 DIN2 N1N258 VDD pch W=1.7U L=0.24U
M4 N1N260 DIN4 N1N268 VDD pch W=1.7U L=0.24U
M3 VDD DIN3 N1N260 VDD pch W=1.8U L=0.24U
M6 N1N278 DIN3 VSS VSS nch W=0.8U L=0.24U
M8 VSS DIN4 N1N278 VSS nch W=0.8U L=0.24U
M7 N1N278 DIN2 N1N268 VSS nch W=0.8U L=0.24U
M10 N1N295 N1N268 VSS VSS nch W=1.2U L=0.24U
M9 N1N295 N1N268 VDD VDD pch W=2.3U L=0.24U
M11 Q N1N295 VDD VDD pch W=4.3U L=0.24U
M12 Q N1N295 VSS VSS nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai24s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N311 VSS nch W=0.8U L=0.24U
M1 N1N301 DIN1 VDD VDD pch W=2.3U L=0.24U
M3 Q DIN2 N1N301 VDD pch W=2.1U L=0.24U
M2 VDD DIN3 N1N303 VDD pch W=4.4U L=0.24U
M4 N1N303 DIN4 N1N305 VDD pch W=4.4U L=0.24U
M5 N1N305 DIN5 N1N307 VDD pch W=4.2U L=0.24U
M6 N1N307 DIN6 Q VDD pch W=4.2U L=0.24U
M9 N1N311 DIN3 VSS VSS nch W=0.8U L=0.24U
M8 N1N311 DIN2 Q VSS nch W=0.8U L=0.24U
M10 VSS DIN6 N1N311 VSS nch W=0.8U L=0.24U
M11 N1N311 DIN4 VSS VSS nch W=0.8U L=0.24U
M12 VSS DIN5 N1N311 VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai24s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N311 VSS nch W=1.3U L=0.24U
M1 N1N301 DIN1 VDD VDD pch W=3.5U L=0.24U
M3 Q DIN2 N1N301 VDD pch W=3.4U L=0.24U
M2 VDD DIN3 N1N303 VDD pch W=6.6U L=0.24U
M4 N1N303 DIN4 N1N305 VDD pch W=6.6U L=0.24U
M5 N1N305 DIN5 N1N307 VDD pch W=6.4U L=0.24U
M6 N1N307 DIN6 Q VDD pch W=6.4U L=0.24U
M9 N1N311 DIN3 VSS VSS nch W=1.3U L=0.24U
M8 N1N311 DIN2 Q VSS nch W=1.3U L=0.24U
M10 VSS DIN6 N1N311 VSS nch W=1.3U L=0.24U
M11 N1N311 DIN4 VSS VSS nch W=1.3U L=0.24U
M12 VSS DIN5 N1N311 VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai24s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N311 VSS nch W=2.14U L=0.24U
M1 N1N301 DIN1 VDD VDD pch W=5.3U L=0.24U
M3 Q DIN2 N1N301 VDD pch W=5.2U L=0.24U
M2 VDD DIN3 N1N303 VDD pch W=9.9U L=0.24U
M4 N1N303 DIN4 N1N305 VDD pch W=9.9U L=0.24U
M5 N1N305 DIN5 N1N307 VDD pch W=9.8U L=0.24U
M6 N1N307 DIN6 Q VDD pch W=9.8U L=0.24U
M9 N1N311 DIN3 VSS VSS nch W=2.14U L=0.24U
M8 N1N311 DIN2 Q VSS nch W=2.14U L=0.24U
M10 VSS DIN6 N1N311 VSS nch W=2.14U L=0.24U
M11 N1N311 DIN4 VSS VSS nch W=2.14U L=0.24U
M12 VSS DIN5 N1N311 VSS nch W=2.14U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai321s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M12 N1N284 DIN3 VSS VSS nch W=1.1U L=0.24U
M6 Q DIN3 N1N257 VDD pch W=2.9U L=0.24U
M5 N1N257 DIN2 N1N256 VDD pch W=3U L=0.24U
M4 N1N256 DIN1 VDD VDD pch W=3.1U L=0.24U
M3 Q DIN6 VDD VDD pch W=1U L=0.24U
M2 Q DIN5 N1N278 VDD pch W=2U L=0.24U
M11 N1N284 DIN1 VSS VSS nch W=1.1U L=0.24U
M9 N1N282 DIN4 N1N284 VSS nch W=1U L=0.24U
M10 N1N284 DIN2 VSS VSS nch W=1.1U L=0.24U
M7 Q DIN6 N1N282 VSS nch W=1U L=0.24U
M8 N1N282 DIN5 N1N284 VSS nch W=1U L=0.24U
M1 N1N278 DIN4 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai321s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M12 N1N284 DIN3 VSS VSS nch W=1.1U L=0.24U
M6 N1N280 DIN3 N1N257 VDD pch W=2.9U L=0.24U
M5 N1N257 DIN2 N1N256 VDD pch W=3U L=0.24U
M4 N1N256 DIN1 VDD VDD pch W=3.1U L=0.24U
M3 N1N280 DIN6 VDD VDD pch W=1U L=0.24U
M2 N1N280 DIN5 N1N278 VDD pch W=2U L=0.24U
M1 N1N278 DIN4 VDD VDD pch W=2U L=0.24U
M11 N1N284 DIN1 VSS VSS nch W=1.1U L=0.24U
M9 N1N282 DIN4 N1N284 VSS nch W=1U L=0.24U
M10 N1N284 DIN2 VSS VSS nch W=1.1U L=0.24U
M7 N1N280 DIN6 N1N282 VSS nch W=1U L=0.24U
M8 N1N282 DIN5 N1N284 VSS nch W=1U L=0.24U
M14 N1N325 N1N280 VSS VSS nch W=0.64U L=0.24U
M13 N1N325 N1N280 VDD VDD pch W=1.4U L=0.24U
M15 Q N1N325 VDD VDD pch W=2.4U L=0.24U
M16 Q N1N325 VSS VSS nch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai321s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M12 N1N284 DIN3 VSS VSS nch W=1.2U L=0.24U
M6 N1N280 DIN3 N1N257 VDD pch W=2.9U L=0.24U
M5 N1N257 DIN2 N1N256 VDD pch W=3U L=0.24U
M4 N1N256 DIN1 VDD VDD pch W=3.1U L=0.24U
M3 N1N280 DIN6 VDD VDD pch W=1U L=0.24U
M2 N1N280 DIN5 N1N278 VDD pch W=2U L=0.24U
M1 N1N278 DIN4 VDD VDD pch W=2U L=0.24U
M11 N1N284 DIN1 VSS VSS nch W=1.2U L=0.24U
M9 N1N282 DIN4 N1N284 VSS nch W=1.1U L=0.24U
M10 N1N284 DIN2 VSS VSS nch W=1.2U L=0.24U
M7 N1N280 DIN6 N1N282 VSS nch W=1U L=0.24U
M8 N1N282 DIN5 N1N284 VSS nch W=1.1U L=0.24U
M14 N1N322 N1N280 VSS VSS nch W=1.1U L=0.24U
M13 N1N322 N1N280 VDD VDD pch W=2.52U L=0.24U
M15 Q N1N322 VDD VDD pch W=4.2U L=0.24U
M16 Q N1N322 VSS VSS nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai322s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M3 Q DIN6 N1N322 VSS nch W=1U L=0.24U
M1 N1N307 DIN4 VDD VDD pch W=1.5U L=0.24U
M2 Q DIN5 N1N307 VDD pch W=1.5U L=0.24U
M6 N1N311 DIN6 VDD VDD pch W=1.5U L=0.24U
M7 Q DIN7 N1N311 VDD pch W=1.5U L=0.24U
M4 N1N322 DIN5 N1N326 VSS nch W=1U L=0.24U
M5 N1N326 DIN2 VSS VSS nch W=1U L=0.24U
M8 Q DIN7 N1N322 VSS nch W=1U L=0.24U
M9 N1N322 DIN4 N1N326 VSS nch W=1U L=0.24U
M10 N1N326 DIN1 VSS VSS nch W=1U L=0.24U
M11 N1N318 DIN1 VDD VDD pch W=2.3U L=0.24U
M12 N1N320 DIN2 N1N318 VDD pch W=2.3U L=0.24U
M13 Q DIN3 N1N320 VDD pch W=2.3U L=0.24U
M14 N1N326 DIN3 VSS VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai322s2 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M3 N1N309 DIN6 N1N322 VSS nch W=1U L=0.24U
M1 N1N307 DIN4 VDD VDD pch W=1.5U L=0.24U
M2 N1N309 DIN5 N1N307 VDD pch W=1.5U L=0.24U
M6 N1N311 DIN6 VDD VDD pch W=1.5U L=0.24U
M7 N1N309 DIN7 N1N311 VDD pch W=1.5U L=0.24U
M4 N1N322 DIN5 N1N326 VSS nch W=1.1U L=0.24U
M5 N1N326 DIN2 VSS VSS nch W=1.1U L=0.24U
M8 N1N309 DIN7 N1N322 VSS nch W=1U L=0.24U
M9 N1N322 DIN4 N1N326 VSS nch W=1.1U L=0.24U
M10 N1N326 DIN1 VSS VSS nch W=1.1U L=0.24U
M11 N1N318 DIN1 VDD VDD pch W=2.3U L=0.24U
M12 N1N320 DIN2 N1N318 VDD pch W=2.3U L=0.24U
M13 N1N309 DIN3 N1N320 VDD pch W=2.3U L=0.24U
M14 N1N326 DIN3 VSS VSS nch W=1.1U L=0.24U
M15 N1N360 N1N309 VDD VDD pch W=2.7U L=0.24U
M16 N1N360 N1N309 VSS VSS nch W=1.1U L=0.24U
M18 Q N1N360 VSS VSS nch W=2.3U L=0.24U
M17 Q N1N360 VDD VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai322s3 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M3 N1N309 DIN6 N1N322 VSS nch W=1.1U L=0.24U
M1 N1N307 DIN4 VDD VDD pch W=1.8U L=0.24U
M2 N1N309 DIN5 N1N307 VDD pch W=1.8U L=0.24U
M6 N1N311 DIN6 VDD VDD pch W=1.8U L=0.24U
M7 N1N309 DIN7 N1N311 VDD pch W=1.8U L=0.24U
M4 N1N322 DIN5 N1N326 VSS nch W=1.3U L=0.24U
M5 N1N326 DIN2 VSS VSS nch W=1.3U L=0.24U
M8 N1N309 DIN7 N1N322 VSS nch W=1.1U L=0.24U
M9 N1N322 DIN4 N1N326 VSS nch W=1.3U L=0.24U
M10 N1N326 DIN1 VSS VSS nch W=1.3U L=0.24U
M11 N1N318 DIN1 VDD VDD pch W=2.7U L=0.24U
M12 N1N320 DIN2 N1N318 VDD pch W=2.7U L=0.24U
M13 N1N309 DIN3 N1N320 VDD pch W=2.7U L=0.24U
M14 N1N326 DIN3 VSS VSS nch W=1.3U L=0.24U
M15 N1N360 N1N309 VDD VDD pch W=4.2U L=0.24U
M16 N1N360 N1N309 VSS VSS nch W=1.7U L=0.24U
M18 Q N1N360 VSS VSS nch W=3.6U L=0.24U
M17 Q N1N360 VDD VDD pch W=6.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai32s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN5 N1N333 VSS nch W=0.8U L=0.24U
M1 N1N321 DIN1 VDD VDD pch W=3.2U L=0.24U
M2 N1N323 DIN2 N1N321 VDD pch W=3.2U L=0.24U
M3 Q DIN3 N1N323 VDD pch W=3.2U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2.1U L=0.24U
M5 N1N327 DIN5 Q VDD pch W=2.1U L=0.24U
M8 N1N333 DIN1 VSS VSS nch W=0.8U L=0.24U
M9 VSS DIN2 N1N333 VSS nch W=0.8U L=0.24U
M7 N1N333 DIN4 Q VSS nch W=0.8U L=0.24U
M10 VSS DIN3 N1N333 VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai32s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN5 N1N333 VSS nch W=1U L=0.24U
M1 N1N321 DIN1 VDD VDD pch W=4.1U L=0.24U
M2 N1N323 DIN2 N1N321 VDD pch W=4U L=0.24U
M3 Q DIN3 N1N323 VDD pch W=3.9U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2.6U L=0.24U
M5 N1N327 DIN5 Q VDD pch W=2.5U L=0.24U
M8 N1N333 DIN1 VSS VSS nch W=1U L=0.24U
M9 VSS DIN2 N1N333 VSS nch W=1U L=0.24U
M7 N1N333 DIN4 Q VSS nch W=1U L=0.24U
M10 VSS DIN3 N1N333 VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai32s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N325 DIN5 N1N333 VSS nch W=0.9U L=0.24U
M1 N1N321 DIN1 VDD VDD pch W=3.1U L=0.24U
M2 N1N323 DIN2 N1N321 VDD pch W=3.1U L=0.24U
M3 N1N325 DIN3 N1N323 VDD pch W=3.1U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2U L=0.24U
M5 N1N327 DIN5 N1N325 VDD pch W=2U L=0.24U
M8 N1N333 DIN1 VSS VSS nch W=0.9U L=0.24U
M9 VSS DIN2 N1N333 VSS nch W=0.9U L=0.24U
M7 N1N333 DIN4 N1N325 VSS nch W=0.9U L=0.24U
M10 VSS DIN3 N1N333 VSS nch W=0.9U L=0.24U
M11 N1N369 N1N325 VDD VDD pch W=2.5U L=0.24U
M13 Q N1N369 VDD VDD pch W=4.5U L=0.24U
M12 N1N369 N1N325 VSS VSS nch W=1.4U L=0.24U
M14 Q N1N369 VSS VSS nch W=2.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai33s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N335 VSS nch W=0.9U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=3.1U L=0.24U
M2 N1N331 DIN2 N1N323 VDD pch W=3U L=0.24U
M3 Q DIN3 N1N331 VDD pch W=2.9U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=3.1U L=0.24U
M5 N1N327 DIN5 N1N329 VDD pch W=3U L=0.24U
M6 N1N329 DIN6 Q VDD pch W=2.9U L=0.24U
M8 N1N335 DIN4 VSS VSS nch W=1.1U L=0.24U
M9 Q DIN2 N1N335 VSS nch W=0.9U L=0.24U
M10 N1N335 DIN5 VSS VSS nch W=1.1U L=0.24U
M11 N1N335 DIN3 Q VSS nch W=0.9U L=0.24U
M12 VSS DIN6 N1N335 VSS nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai33s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N333 DIN1 N1N335 VSS nch W=0.8U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N331 DIN2 N1N323 VDD pch W=1.9U L=0.24U
M3 N1N333 DIN3 N1N331 VDD pch W=1.9U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2.1U L=0.24U
M5 N1N327 DIN5 N1N329 VDD pch W=1.9U L=0.24U
M6 N1N329 DIN6 N1N333 VDD pch W=1.9U L=0.24U
M8 N1N335 DIN4 VSS VSS nch W=0.9U L=0.24U
M9 N1N333 DIN2 N1N335 VSS nch W=0.8U L=0.24U
M10 N1N335 DIN5 VSS VSS nch W=0.9U L=0.24U
M11 N1N335 DIN3 N1N333 VSS nch W=0.8U L=0.24U
M12 VSS DIN6 N1N335 VSS nch W=0.9U L=0.24U
M13 N1N383 N1N333 VDD VDD pch W=1.1U L=0.24U
M14 N1N383 N1N333 VSS VSS nch W=0.6U L=0.24U
M15 Q N1N383 VDD VDD pch W=2.4U L=0.24U
M16 Q N1N383 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT oai33s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N333 DIN1 N1N335 VSS nch W=0.8U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N331 DIN2 N1N323 VDD pch W=1.9U L=0.24U
M3 N1N333 DIN3 N1N331 VDD pch W=1.9U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2.1U L=0.24U
M5 N1N327 DIN5 N1N329 VDD pch W=1.9U L=0.24U
M6 N1N329 DIN6 N1N333 VDD pch W=1.9U L=0.24U
M8 N1N335 DIN4 VSS VSS nch W=0.9U L=0.24U
M9 N1N333 DIN2 N1N335 VSS nch W=0.8U L=0.24U
M10 N1N335 DIN5 VSS VSS nch W=0.9U L=0.24U
M11 N1N335 DIN3 N1N333 VSS nch W=0.8U L=0.24U
M12 VSS DIN6 N1N335 VSS nch W=0.9U L=0.24U
M13 N1N383 N1N333 VDD VDD pch W=2U L=0.24U
M14 N1N383 N1N333 VSS VSS nch W=1U L=0.24U
M15 Q N1N383 VDD VDD pch W=4.2U L=0.24U
M16 Q N1N383 VSS VSS nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or2s1 Q DIN1 DIN2
M3 N1N441 DIN1 VSS VSS nch W=0.7U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=1.6U L=0.24U
M2 N1N441 DIN2 N1N428 VDD pch W=1.6U L=0.24U
M4 N1N441 DIN2 VSS VSS nch W=0.7U L=0.24U
M6 Q N1N441 VSS VSS nch W=1.3U L=0.24U
M5 Q N1N441 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or2s2 Q DIN1 DIN2
M3 N1N441 DIN1 VSS VSS nch W=1.1U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=3U L=0.24U
M2 N1N441 DIN2 N1N428 VDD pch W=3U L=0.24U
M4 N1N441 DIN2 VSS VSS nch W=1.1U L=0.24U
M6 Q N1N441 VSS VSS nch W=3.5U L=0.24U
M5 Q N1N441 VDD VDD pch W=4.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or2s3 Q DIN1 DIN2
M3 N1N441 DIN1 VSS VSS nch W=2.2U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=5.8U L=0.24U
M2 N1N441 DIN2 N1N428 VDD pch W=5.8U L=0.24U
M4 N1N441 DIN2 VSS VSS nch W=2.2U L=0.24U
M6 Q N1N441 VSS VSS nch W=6.2U L=0.24U
M5 Q N1N441 VDD VDD pch W=7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or3s1 Q DIN1 DIN2 DIN3
M4 N1N434 DIN1 VSS VSS nch W=0.7U L=0.24U
M1 N1N430 DIN1 VDD VDD pch W=3.16U L=0.24U
M2 N1N432 DIN2 N1N430 VDD pch W=3.16U L=0.24U
M3 N1N434 DIN3 N1N432 VDD pch W=3.16U L=0.24U
M5 N1N434 DIN2 VSS VSS nch W=0.7U L=0.24U
M6 N1N434 DIN3 VSS VSS nch W=0.7U L=0.24U
M7 Q N1N434 VDD VDD pch W=2.1U L=0.24U
M8 Q N1N434 VSS VSS nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or3s2 Q DIN1 DIN2 DIN3
M4 N1N434 DIN1 VSS VSS nch W=1.1U L=0.24U
M1 N1N430 DIN1 VDD VDD pch W=4.2U L=0.24U
M2 N1N432 DIN2 N1N430 VDD pch W=4.1U L=0.24U
M3 N1N434 DIN3 N1N432 VDD pch W=4U L=0.24U
M5 N1N434 DIN2 VSS VSS nch W=1.1U L=0.24U
M6 N1N434 DIN3 VSS VSS nch W=1.1U L=0.24U
M7 Q N1N434 VDD VDD pch W=5.2U L=0.24U
M8 Q N1N434 VSS VSS nch W=4.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or3s3 Q DIN1 DIN2 DIN3
M4 N1N434 DIN1 VSS VSS nch W=2U L=0.24U
M1 N1N430 DIN1 VDD VDD pch W=8.5U L=0.24U
M2 N1N432 DIN2 N1N430 VDD pch W=7.8U L=0.24U
M3 N1N434 DIN3 N1N432 VDD pch W=6.2U L=0.24U
M5 N1N434 DIN2 VSS VSS nch W=2U L=0.24U
M6 N1N434 DIN3 VSS VSS nch W=2U L=0.24U
M7 Q N1N434 VDD VDD pch W=7.1U L=0.24U
M8 Q N1N434 VSS VSS nch W=6.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or4s1 Q DIN1 DIN2 DIN3 DIN4
M5 N1N438 DIN1 VSS VSS nch W=0.7U L=0.24U
M1 N1N432 DIN1 VDD VDD pch W=4.5U L=0.24U
M2 N1N434 DIN2 N1N432 VDD pch W=4.2U L=0.24U
M3 N1N436 DIN3 N1N434 VDD pch W=4.1U L=0.24U
M4 N1N438 DIN4 N1N436 VDD pch W=3.1U L=0.24U
M6 N1N438 DIN2 VSS VSS nch W=0.7U L=0.24U
M7 N1N438 DIN3 VSS VSS nch W=0.7U L=0.24U
M8 N1N438 DIN4 VSS VSS nch W=0.7U L=0.24U
M9 Q N1N438 VDD VDD pch W=2.3U L=0.24U
M10 Q N1N438 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or4s2 Q DIN1 DIN2 DIN3 DIN4
M5 N1N438 DIN1 VSS VSS nch W=1.56U L=0.24U
M1 N1N432 DIN1 VDD VDD pch W=9.5U L=0.24U
M2 N1N434 DIN2 N1N432 VDD pch W=9.2U L=0.24U
M3 N1N436 DIN3 N1N434 VDD pch W=9U L=0.24U
M4 N1N438 DIN4 N1N436 VDD pch W=8.5U L=0.24U
M6 N1N438 DIN2 VSS VSS nch W=1.56U L=0.24U
M7 N1N438 DIN3 VSS VSS nch W=1.56U L=0.24U
M8 N1N438 DIN4 VSS VSS nch W=1.56U L=0.24U
M9 Q N1N438 VDD VDD pch W=6.3U L=0.24U
M10 Q N1N438 VSS VSS nch W=3.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or4s3 Q DIN1 DIN2 DIN3 DIN4
M1 N1N425 DIN1 VDD VDD pch W=4.4U L=0.24U
M2 N1N441 DIN2 N1N425 VDD pch W=3.9U L=0.24U
M3 N1N441 DIN1 VSS VSS nch W=1.7U L=0.24U
M4 N1N441 DIN2 VSS VSS nch W=1.7U L=0.24U
M5 N1N422 DIN3 VDD VDD pch W=4.4U L=0.24U
M6 N1N428 DIN4 N1N422 VDD pch W=3.9U L=0.24U
M7 N1N428 DIN3 VSS VSS nch W=1.7U L=0.24U
M8 N1N428 DIN4 VSS VSS nch W=1.7U L=0.24U
M9 Q N1N441 VDD VDD pch W=4.2U L=0.24U
M11 Q N1N441 N1N445 VSS nch W=4.2U L=0.24U
M12 N1N445 N1N428 VSS VSS nch W=4.2U L=0.24U
M10 VDD N1N428 Q VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or5s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 VSS VSS nch W=0.7U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=3U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=2.6U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=2.4U L=0.24U
M4 N1N444 DIN3 VSS VSS nch W=0.7U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=0.7U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=1.9U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=1.7U L=0.24U
M9 N1N494 DIN5 VSS VSS nch W=0.7U L=0.24U
M10 VSS DIN4 N1N494 VSS nch W=0.7U L=0.24U
M11 Q N1N444 VDD VDD pch W=2U L=0.24U
M12 VDD N1N494 Q VDD pch W=2U L=0.24U
M13 Q N1N444 N1N480 VSS nch W=1.7U L=0.24U
M14 N1N480 N1N494 VSS VSS nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or5s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 VSS VSS nch W=1.4U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=6U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=5.8U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=5.6U L=0.24U
M4 N1N444 DIN3 VSS VSS nch W=1.4U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=1.4U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=3.9U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=3.7U L=0.24U
M9 N1N494 DIN5 VSS VSS nch W=1.4U L=0.24U
M10 VSS DIN4 N1N494 VSS nch W=1.4U L=0.24U
M11 Q N1N444 VDD VDD pch W=4U L=0.24U
M12 VDD N1N494 Q VDD pch W=4U L=0.24U
M13 Q N1N444 N1N480 VSS nch W=3.6U L=0.24U
M14 N1N480 N1N494 VSS VSS nch W=3.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT or5s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 VSS VSS nch W=2.3U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=10.6U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=9.9U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=9.4U L=0.24U
M4 N1N444 DIN3 VSS VSS nch W=2.3U L=0.24U
M6 N1N444 DIN1 VSS VSS nch W=2.3U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=6.34U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=6.2U L=0.24U
M9 N1N494 DIN5 VSS VSS nch W=2.3U L=0.24U
M10 VSS DIN4 N1N494 VSS nch W=2.3U L=0.24U
M11 Q N1N444 VDD VDD pch W=6.8U L=0.24U
M12 VDD N1N494 Q VDD pch W=6.8U L=0.24U
M13 Q N1N444 N1N480 VSS nch W=5.7U L=0.24U
M14 N1N480 N1N494 VSS VSS nch W=5.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ppt1s1 OUTD DIN OUTS
M1 OUTD DIN OUTS VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ppt1s2 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ppt1s3 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ppt1s4 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ppt1s5 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=32U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ppt1s6 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ppu1s1 OUTD GIN
M1 OUTD GIN VDD VDD pch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ppu1s2 OUTD GIN
M1 OUTD GIN VDD VDD pch W=3.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT rpc1s1 DIN
M1 N1N254 N1N294 VDD VDD pch W=0.8U L=0.24U
M3 DIN N1N294 N1N258 VSS nch W=0.8U L=0.24U
M2 DIN N1N294 N1N254 VDD pch W=0.8U L=0.24U
M4 N1N258 N1N294 VSS VSS nch W=0.8U L=0.24U
M5 N1N294 DIN VDD VDD pch W=1.6U L=0.24U
M6 N1N294 DIN VSS VSS nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT rpc1s2 DIN
M1 N1N254 N1N294 VDD VDD pch W=1.2U L=0.24U
M3 DIN N1N294 N1N258 VSS nch W=1.2U L=0.24U
M2 DIN N1N294 N1N254 VDD pch W=1.2U L=0.24U
M4 N1N258 N1N294 VSS VSS nch W=1.2U L=0.24U
M5 N1N294 DIN VDD VDD pch W=2.5U L=0.24U
M6 N1N294 DIN VSS VSS nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffacs1 Q QN CLRB CLK SSEL SDIN DIN
M23 TP7 CLRB VDD VDD pch W=1.3U L=0.24U
M27 Q TP8 VDD VDD pch W=3.14U L=0.24U
M15 TP5 TP3 VDD VDD pch W=1.3U L=0.24U
M30 QN Q VSS VSS nch W=1.42U L=0.24U
M9 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M10 TP21 TP1 TP3 VSS nch W=0.8U L=0.24U
M19 TP5 CLK TP8 VSS nch W=0.96U L=0.24U
M20 TP8 TP1 TP5 VDD pch W=1.4U L=0.24U
M12 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M21 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M22 TP8 TP1 TP7 VSS nch W=0.8U L=0.24U
M29 QN Q VDD VDD pch W=3.02U L=0.24U
M11 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M17 TP5 TP3 TP6 VSS nch W=0.9U L=0.24U
M25 TP7 Q TP9 VSS nch W=0.9U L=0.24U
M28 Q TP8 VSS VSS nch W=1.96U L=0.24U
M16 TP5 CLRB VDD VDD pch W=1.3U L=0.24U
M14 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M18 TP6 CLRB VSS VSS nch W=0.9U L=0.24U
M7 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M24 TP7 Q VDD VDD pch W=1.3U L=0.24U
M26 TP9 CLRB VSS VSS nch W=0.9U L=0.24U
M8 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffacs2 Q QN CLRB CLK SSEL SDIN DIN
M23 TP7 CLRB VDD VDD pch W=1.3U L=0.24U
M27 Q TP8 VDD VDD pch W=6.2U L=0.24U
M15 TP5 TP3 VDD VDD pch W=1.84U L=0.24U
M30 QN Q VSS VSS nch W=2.68U L=0.24U
M9 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M10 TP21 TP1 TP3 VSS nch W=0.8U L=0.24U
M19 TP5 CLK TP8 VSS nch W=1.52U L=0.24U
M20 TP8 TP1 TP5 VDD pch W=1.9U L=0.24U
M12 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M21 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M22 TP8 TP1 TP7 VSS nch W=0.8U L=0.24U
M29 QN Q VDD VDD pch W=6.16U L=0.24U
M11 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M17 TP5 TP3 TP6 VSS nch W=1.48U L=0.24U
M25 TP7 Q TP9 VSS nch W=0.9U L=0.24U
M28 Q TP8 VSS VSS nch W=3.98U L=0.24U
M16 TP5 CLRB VDD VDD pch W=1.84U L=0.24U
M14 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M18 TP6 CLRB VSS VSS nch W=1.48U L=0.24U
M7 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M24 TP7 Q VDD VDD pch W=1.3U L=0.24U
M26 TP9 CLRB VSS VSS nch W=0.9U L=0.24U
M8 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffascs1 SETB CLRB DIN SSEL SDIN CLK QN Q
M18 TP6 CLK VSS VSS nch W=0.8U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M12 TP0 SETB VSS VSS nch W=0.8U L=0.24U
M8 TP1 CLRB VSS VSS nch W=0.8U L=0.24U
M7 TP1 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP1 VDD VDD pch W=2.2U L=0.24U
M10 TP4 TP1 VSS VSS nch W=1.4U L=0.24U
M39 Q TP13 VDD VDD pch W=3.18U L=0.24U
M29 TP11 TP8 TP12 VSS nch W=2.2U L=0.24U
M19 TP8 CLK TP21 VDD pch W=1.3U L=0.24U
M20 TP21 TP6 TP8 VSS nch W=0.8U L=0.24U
M31 TP11 CLK TP13 VSS nch W=2.2U L=0.24U
M32 TP13 TP6 TP11 VDD pch W=2.5U L=0.24U
M21 TP8 CLK TP9 VSS nch W=0.8U L=0.24U
M22 TP9 TP6 TP8 VDD pch W=1.3U L=0.24U
M33 TP14 CLK TP13 VDD pch W=1.3U L=0.24U
M27 TP11 TP8 VDD VDD pch W=2.4U L=0.24U
M28 TP11 TP4 VDD VDD pch W=2.4U L=0.24U
M26 TP10 TP11 VSS VSS nch W=0.8U L=0.24U
M38 TP15 TP4 VSS VSS nch W=0.8U L=0.24U
M30 TP12 TP4 VSS VSS nch W=2.2U L=0.24U
M42 TP16 TP13 VSS VSS nch W=2.64U L=0.24U
M40 Q TP2 VDD VDD pch W=3.18U L=0.24U
M41 Q TP2 TP16 VSS nch W=2.64U L=0.24U
M25 TP9 TP2 TP10 VSS nch W=0.8U L=0.24U
M17 TP6 CLK VDD VDD pch W=1.4U L=0.24U
M15 TP2 TP0 TP3 VSS nch W=1.3U L=0.24U
M16 TP3 TP4 VSS VSS nch W=1.3U L=0.24U
M44 QN Q VSS VSS nch W=1.44U L=0.24U
M13 TP2 TP0 VDD VDD pch W=1.8U L=0.24U
M14 TP2 TP4 VDD VDD pch W=1.8U L=0.24U
M23 TP9 TP2 VDD VDD pch W=1.3U L=0.24U
M24 TP9 TP11 VDD VDD pch W=1.3U L=0.24U
M37 TP14 Q TP15 VSS nch W=0.8U L=0.24U
M36 TP14 Q VDD VDD pch W=1.3U L=0.24U
M34 TP13 TP6 TP14 VSS nch W=0.8U L=0.24U
M43 QN Q VDD VDD pch W=3.18U L=0.24U
M11 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M35 TP14 TP4 VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffascs2 SETB CLRB DIN SSEL SDIN CLK QN Q
M18 TP6 CLK VSS VSS nch W=0.8U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M12 TP0 SETB VSS VSS nch W=0.8U L=0.24U
M8 TP1 CLRB VSS VSS nch W=0.8U L=0.24U
M7 TP1 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP1 VDD VDD pch W=2.7U L=0.24U
M10 TP4 TP1 VSS VSS nch W=2.2U L=0.24U
M39 Q TP13 VDD VDD pch W=6.26U L=0.24U
M29 TP11 TP8 TP12 VSS nch W=2.92U L=0.24U
M19 TP8 CLK TP21 VDD pch W=1.3U L=0.24U
M20 TP21 TP6 TP8 VSS nch W=0.8U L=0.24U
M31 TP11 CLK TP13 VSS nch W=2.7U L=0.24U
M32 TP13 TP6 TP11 VDD pch W=3U L=0.24U
M21 TP8 CLK TP9 VSS nch W=0.8U L=0.24U
M22 TP9 TP6 TP8 VDD pch W=1.3U L=0.24U
M33 TP14 CLK TP13 VDD pch W=1.3U L=0.24U
M27 TP11 TP8 VDD VDD pch W=3.24U L=0.24U
M28 TP11 TP4 VDD VDD pch W=3.24U L=0.24U
M26 TP10 TP11 VSS VSS nch W=0.8U L=0.24U
M38 TP15 TP4 VSS VSS nch W=0.8U L=0.24U
M30 TP12 TP4 VSS VSS nch W=2.92U L=0.24U
M42 TP16 TP13 VSS VSS nch W=5.26U L=0.24U
M40 Q TP2 VDD VDD pch W=6.26U L=0.24U
M41 Q TP2 TP16 VSS nch W=5.26U L=0.24U
M25 TP9 TP2 TP10 VSS nch W=0.8U L=0.24U
M17 TP6 CLK VDD VDD pch W=1.6U L=0.24U
M15 TP2 TP0 TP3 VSS nch W=2.2U L=0.24U
M16 TP3 TP4 VSS VSS nch W=2.2U L=0.24U
M44 QN Q VSS VSS nch W=2.88U L=0.24U
M13 TP2 TP0 VDD VDD pch W=2.82U L=0.24U
M14 TP2 TP4 VDD VDD pch W=2.82U L=0.24U
M23 TP9 TP2 VDD VDD pch W=1.3U L=0.24U
M24 TP9 TP11 VDD VDD pch W=1.3U L=0.24U
M37 TP14 Q TP15 VSS nch W=0.8U L=0.24U
M36 TP14 Q VDD VDD pch W=1.3U L=0.24U
M34 TP13 TP6 TP14 VSS nch W=0.8U L=0.24U
M43 QN Q VDD VDD pch W=6.2U L=0.24U
M11 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M35 TP14 TP4 VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffass1 Q QN SETB CLK SSEL SDIN DIN
M27 TP7 SETB VDD VDD pch W=1.3U L=0.24U
M19 TP5 TP3 VDD VDD pch W=1.3U L=0.24U
M34 Q QN VSS VSS nch W=1.42U L=0.24U
M13 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M14 TP21 TP1 TP3 VSS nch W=0.8U L=0.24U
M23 TP5 CLK TP8 VSS nch W=0.96U L=0.24U
M24 TP8 TP1 TP5 VDD pch W=1.4U L=0.24U
M16 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M25 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M33 Q QN VDD VDD pch W=3.02U L=0.24U
M15 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M29 TP7 QN TP9 VSS nch W=0.9U L=0.24U
M32 QN TP8 VSS VSS nch W=1.96U L=0.24U
M20 TP5 SETB VDD VDD pch W=1.3U L=0.24U
M18 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M22 TP6 SETB VSS VSS nch W=0.9U L=0.24U
M17 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M30 TP9 SETB VSS VSS nch W=0.9U L=0.24U
M28 TP7 QN VDD VDD pch W=1.3U L=0.24U
M21 TP5 TP3 TP6 VSS nch W=0.9U L=0.24U
M12 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M26 TP8 TP1 TP7 VSS nch W=0.8U L=0.24U
M31 QN TP8 VDD VDD pch W=3.14U L=0.24U
M11 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M3 TP19 SDIN VDD VDD pch W=1.3U L=0.24U
M4 TP19 SDIN VSS VSS nch W=0.8U L=0.24U
M1 TP18 DIN VDD VDD pch W=1.3U L=0.24U
M2 TP18 DIN VSS VSS nch W=0.8U L=0.24U
M9 TP21 TP20 TP19 VDD pch W=1.3U L=0.24U
M10 TP19 SSEL TP21 VSS nch W=0.8U L=0.24U
M5 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M6 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M8 TP18 TP20 TP21 VSS nch W=0.8U L=0.24U
M7 TP21 SSEL TP18 VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffass2 Q QN SETB CLK SSEL SDIN DIN
M27 TP7 SETB VDD VDD pch W=1.3U L=0.24U
M19 TP5 TP3 VDD VDD pch W=1.84U L=0.24U
M34 Q QN VSS VSS nch W=2.68U L=0.24U
M13 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M14 TP21 TP1 TP3 VSS nch W=0.8U L=0.24U
M23 TP5 CLK TP8 VSS nch W=1.52U L=0.24U
M24 TP8 TP1 TP5 VDD pch W=1.9U L=0.24U
M16 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M25 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M33 Q QN VDD VDD pch W=6.16U L=0.24U
M15 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M29 TP7 QN TP9 VSS nch W=0.9U L=0.24U
M32 QN TP8 VSS VSS nch W=3.98U L=0.24U
M20 TP5 SETB VDD VDD pch W=1.84U L=0.24U
M18 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M22 TP6 SETB VSS VSS nch W=1.48U L=0.24U
M17 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M30 TP9 SETB VSS VSS nch W=0.9U L=0.24U
M28 TP7 QN VDD VDD pch W=1.3U L=0.24U
M21 TP5 TP3 TP6 VSS nch W=1.48U L=0.24U
M12 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M26 TP8 TP1 TP7 VSS nch W=0.8U L=0.24U
M31 QN TP8 VDD VDD pch W=6.2U L=0.24U
M11 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M3 TP19 SDIN VDD VDD pch W=1.3U L=0.24U
M4 TP19 SDIN VSS VSS nch W=0.8U L=0.24U
M1 TP18 DIN VDD VDD pch W=1.3U L=0.24U
M2 TP18 DIN VSS VSS nch W=0.8U L=0.24U
M9 TP21 TP20 TP19 VDD pch W=1.3U L=0.24U
M10 TP19 SSEL TP21 VSS nch W=0.8U L=0.24U
M5 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M6 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M8 TP18 TP20 TP21 VSS nch W=0.8U L=0.24U
M7 TP21 SSEL TP18 VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffcs1 SSEL CLRB DIN SDIN CLK Q QN
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M9 TP2 TP21 TP1 VSS nch W=0.8U L=0.24U
M8 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M7 TP2 TP21 VDD VDD pch W=1.3U L=0.24U
M12 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M13 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M14 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M19 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M21 TP6 CLK TP7 VSS nch W=0.8U L=0.24U
M22 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M27 QN TP7 VDD VDD pch W=3.14U L=0.24U
M28 QN TP7 VSS VSS nch W=2.06U L=0.24U
M15 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M16 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M18 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M23 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M29 Q QN VDD VDD pch W=2.94U L=0.24U
M30 Q QN VSS VSS nch W=1.28U L=0.24U
M20 TP6 TP4 VSS VSS nch W=0.8U L=0.24U
M11 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M26 TP8 QN VSS VSS nch W=0.8U L=0.24U
M24 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M25 TP8 QN VDD VDD pch W=1.3U L=0.24U
M17 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M10 TP1 CLRB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffcs2 SSEL CLRB DIN SDIN CLK Q QN
M13 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M14 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M19 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M21 TP6 CLK TP7 VSS nch W=1.3U L=0.24U
M22 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M27 QN TP7 VDD VDD pch W=6.24U L=0.24U
M28 QN TP7 VSS VSS nch W=3.98U L=0.24U
M15 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M16 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M17 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M18 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M23 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M24 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M25 TP8 QN VDD VDD pch W=1.3U L=0.24U
M26 TP8 QN VSS VSS nch W=0.8U L=0.24U
M29 Q QN VDD VDD pch W=5.92U L=0.24U
M30 Q QN VSS VSS nch W=2.66U L=0.24U
M20 TP6 TP4 VSS VSS nch W=1.26U L=0.24U
M11 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M12 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M7 TP2 TP21 VDD VDD pch W=1.3U L=0.24U
M8 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP2 TP21 TP1 VSS nch W=0.8U L=0.24U
M10 TP1 CLRB VSS VSS nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffles1 EB DIN SSEL SDIN CLK QN Q
M29 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M30 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M40 TP9 TP10 VSS VSS nch W=0.8U L=0.24U
M50 Q TP11 VSS VSS nch W=2.06U L=0.24U
M42 TP10 TP8 VSS VSS nch W=0.8U L=0.24U
M48 TP5 Q VSS VSS nch W=0.8U L=0.24U
M47 TP5 Q VDD VDD pch W=1.3U L=0.24U
M52 QN Q VSS VSS nch W=1.28U L=0.24U
M35 TP8 CLK TP3 VDD pch W=1.3U L=0.24U
M36 TP3 TP7 TP8 VSS nch W=0.8U L=0.24U
M43 TP10 CLK TP11 VSS nch W=0.8U L=0.24U
M38 TP9 TP7 TP8 VDD pch W=1.3U L=0.24U
M46 TP11 TP7 TP5 VSS nch W=0.8U L=0.24U
M51 QN Q VDD VDD pch W=2.94U L=0.24U
M37 TP8 CLK TP9 VSS nch W=0.8U L=0.24U
M49 Q TP11 VDD VDD pch W=3.14U L=0.24U
M41 TP10 TP8 VDD VDD pch W=1.8U L=0.24U
M39 TP9 TP10 VDD VDD pch W=1.3U L=0.24U
M44 TP11 TP7 TP10 VDD pch W=1.3U L=0.24U
M45 TP5 CLK TP11 VDD pch W=1.3U L=0.24U
M19 TP3 TP23 SDIN VDD pch W=1.3U L=0.24U
M20 SDIN SSEL TP3 VSS nch W=0.8U L=0.24U
M28 TP27 TP25 VSS VSS nch W=0.8U L=0.24U
M27 TP27 TP25 VDD VDD pch W=1.3U L=0.24U
M21 TP25 EB VDD VDD pch W=1.3U L=0.24U
M23 TP25 EB TP26 VSS nch W=0.8U L=0.24U
M24 TP26 TP23 VSS VSS nch W=0.8U L=0.24U
M6 TP22 TP23 VSS VSS nch W=0.8U L=0.24U
M18 TP24 TP21 VSS VSS nch W=0.8U L=0.24U
M17 TP24 TP21 VDD VDD pch W=1.3U L=0.24U
M3 TP21 TP20 VDD VDD pch W=1.3U L=0.24U
M5 TP21 TP20 TP22 VSS nch W=0.8U L=0.24U
M2 TP20 EB VSS VSS nch W=0.8U L=0.24U
M1 TP20 EB VDD VDD pch W=1.3U L=0.24U
M15 TP3 TP21 DIN VDD pch W=1.3U L=0.24U
M16 DIN TP24 TP3 VSS nch W=0.8U L=0.24U
M25 TP4 TP25 TP3 VDD pch W=1.3U L=0.24U
M26 TP3 TP27 TP4 VSS nch W=0.8U L=0.24U
M4 TP21 TP23 VDD VDD pch W=1.3U L=0.24U
M22 TP25 TP23 VDD VDD pch W=1.3U L=0.24U
M34 TP7 CLK VSS VSS nch W=0.8U L=0.24U
M33 TP7 CLK VDD VDD pch W=1.3U L=0.24U
M11 TP23 SSEL VDD VDD pch W=1.5U L=0.24U
M12 TP23 SSEL VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffles2 EB DIN SSEL SDIN CLK QN Q
M29 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M30 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M40 TP9 TP10 VSS VSS nch W=0.8U L=0.24U
M50 Q TP11 VSS VSS nch W=3.98U L=0.24U
M42 TP10 TP8 VSS VSS nch W=1.26U L=0.24U
M48 TP5 Q VSS VSS nch W=0.8U L=0.24U
M47 TP5 Q VDD VDD pch W=1.3U L=0.24U
M52 QN Q VSS VSS nch W=2.66U L=0.24U
M35 TP8 CLK TP3 VDD pch W=1.3U L=0.24U
M36 TP3 TP7 TP8 VSS nch W=0.8U L=0.24U
M43 TP10 CLK TP11 VSS nch W=1.3U L=0.24U
M38 TP9 TP7 TP8 VDD pch W=1.3U L=0.24U
M46 TP11 TP7 TP5 VSS nch W=0.8U L=0.24U
M51 QN Q VDD VDD pch W=5.92U L=0.24U
M37 TP8 CLK TP9 VSS nch W=0.8U L=0.24U
M49 Q TP11 VDD VDD pch W=6.24U L=0.24U
M41 TP10 TP8 VDD VDD pch W=2.78U L=0.24U
M39 TP9 TP10 VDD VDD pch W=1.3U L=0.24U
M44 TP11 TP7 TP10 VDD pch W=1.8U L=0.24U
M45 TP5 CLK TP11 VDD pch W=1.3U L=0.24U
M19 TP3 TP23 SDIN VDD pch W=1.3U L=0.24U
M20 SDIN SSEL TP3 VSS nch W=0.8U L=0.24U
M28 TP27 TP25 VSS VSS nch W=0.8U L=0.24U
M27 TP27 TP25 VDD VDD pch W=1.3U L=0.24U
M21 TP25 EB VDD VDD pch W=1.3U L=0.24U
M23 TP25 EB TP26 VSS nch W=0.8U L=0.24U
M24 TP26 TP23 VSS VSS nch W=0.8U L=0.24U
M6 TP22 TP23 VSS VSS nch W=0.8U L=0.24U
M18 TP24 TP21 VSS VSS nch W=0.8U L=0.24U
M17 TP24 TP21 VDD VDD pch W=1.3U L=0.24U
M3 TP21 TP20 VDD VDD pch W=1.3U L=0.24U
M5 TP21 TP20 TP22 VSS nch W=0.8U L=0.24U
M2 TP20 EB VSS VSS nch W=0.8U L=0.24U
M1 TP20 EB VDD VDD pch W=1.3U L=0.24U
M15 TP3 TP21 DIN VDD pch W=1.3U L=0.24U
M16 DIN TP24 TP3 VSS nch W=0.8U L=0.24U
M25 TP4 TP25 TP3 VDD pch W=1.3U L=0.24U
M26 TP3 TP27 TP4 VSS nch W=0.8U L=0.24U
M4 TP21 TP23 VDD VDD pch W=1.3U L=0.24U
M22 TP25 TP23 VDD VDD pch W=1.3U L=0.24U
M34 TP7 CLK VSS VSS nch W=0.8U L=0.24U
M33 TP7 CLK VDD VDD pch W=1.3U L=0.24U
M11 TP23 SSEL VDD VDD pch W=1.5U L=0.24U
M12 TP23 SSEL VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffs1 Q QN CLK SSEL SDIN DIN
M17 TP3 CLK TP9 VDD pch W=1.3U L=0.24U
M18 TP9 TP1 TP3 VSS nch W=0.8U L=0.24U
M21 TP5 TP3 VDD VDD pch W=1.8U L=0.24U
M25 TP5 CLK TP6 VSS nch W=0.8U L=0.24U
M26 TP6 TP1 TP5 VDD pch W=1.3U L=0.24U
M29 Q TP6 VDD VDD pch W=3.14U L=0.24U
M30 Q TP6 VSS VSS nch W=2.06U L=0.24U
M19 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M20 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M23 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M24 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M27 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M28 TP6 TP1 TP7 VSS nch W=0.8U L=0.24U
M31 TP7 Q VDD VDD pch W=1.3U L=0.24U
M32 TP7 Q VSS VSS nch W=0.8U L=0.24U
M33 QN Q VDD VDD pch W=2.94U L=0.24U
M34 QN Q VSS VSS nch W=1.28U L=0.24U
M22 TP5 TP3 VSS VSS nch W=0.8U L=0.24U
M14 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M13 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M9 DIN TP8 TP9 VSS nch W=0.8U L=0.24U
M10 TP9 SSEL DIN VDD pch W=1.3U L=0.24U
M11 TP9 TP8 SDIN VDD pch W=1.3U L=0.24U
M12 SDIN SSEL TP9 VSS nch W=0.8U L=0.24U
M6 TP8 SSEL VSS VSS nch W=0.8U L=0.24U
M5 TP8 SSEL VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffs2 Q QN CLK SSEL SDIN DIN
M17 TP3 CLK TP9 VDD pch W=1.3U L=0.24U
M18 TP9 TP1 TP3 VSS nch W=0.8U L=0.24U
M21 TP5 TP3 VDD VDD pch W=2.76U L=0.24U
M25 TP5 CLK TP6 VSS nch W=1.3U L=0.24U
M26 TP6 TP1 TP5 VDD pch W=1.8U L=0.24U
M29 Q TP6 VDD VDD pch W=6.24U L=0.24U
M30 Q TP6 VSS VSS nch W=3.98U L=0.24U
M19 TP3 CLK TP4 VSS nch W=0.8U L=0.24U
M20 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M23 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M24 TP4 TP5 VSS VSS nch W=0.8U L=0.24U
M27 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M28 TP6 TP1 TP7 VSS nch W=0.8U L=0.24U
M31 TP7 Q VDD VDD pch W=1.3U L=0.24U
M32 TP7 Q VSS VSS nch W=0.8U L=0.24U
M33 QN Q VDD VDD pch W=5.92U L=0.24U
M34 QN Q VSS VSS nch W=2.66U L=0.24U
M22 TP5 TP3 VSS VSS nch W=1.26U L=0.24U
M14 TP1 CLK VSS VSS nch W=0.8U L=0.24U
M13 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M9 DIN TP8 TP9 VSS nch W=0.8U L=0.24U
M10 TP9 SSEL DIN VDD pch W=1.3U L=0.24U
M11 TP9 TP8 SDIN VDD pch W=1.3U L=0.24U
M12 SDIN SSEL TP9 VSS nch W=0.8U L=0.24U
M6 TP8 SSEL VSS VSS nch W=0.8U L=0.24U
M5 TP8 SSEL VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffscs1 SSEL CLR DIN SET SDIN CLK QN Q
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M17 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M18 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M23 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M25 TP6 CLK TP7 VSS nch W=0.8U L=0.24U
M26 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M31 QN TP7 VDD VDD pch W=3.14U L=0.24U
M32 QN TP7 VSS VSS nch W=2.06U L=0.24U
M19 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M20 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M22 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M27 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M33 Q QN VDD VDD pch W=2.94U L=0.24U
M34 Q QN VSS VSS nch W=1.28U L=0.24U
M24 TP6 TP4 VSS VSS nch W=0.8U L=0.24U
M15 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M16 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M30 TP8 QN VSS VSS nch W=0.8U L=0.24U
M28 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M29 TP8 QN VDD VDD pch W=1.3U L=0.24U
M21 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M9 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M10 TP2 TP21 TP1 VDD pch W=1.3U L=0.24U
M11 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M12 TP2 CLRB TP9 VSS nch W=0.8U L=0.24U
M13 TP9 TP21 VSS VSS nch W=0.8U L=0.24U
M14 TP9 TP0 VSS VSS nch W=0.8U L=0.24U
M7 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M8 TP0 SETB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffscs2 SSEL CLR DIN SET SDIN CLK QN Q
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M17 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M18 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M23 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M25 TP6 CLK TP7 VSS nch W=1.3U L=0.24U
M26 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M31 QN TP7 VDD VDD pch W=6.24U L=0.24U
M32 QN TP7 VSS VSS nch W=3.98U L=0.24U
M19 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M20 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M22 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M27 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M33 Q QN VDD VDD pch W=5.92U L=0.24U
M34 Q QN VSS VSS nch W=2.66U L=0.24U
M24 TP6 TP4 VSS VSS nch W=1.26U L=0.24U
M15 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M16 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M30 TP8 QN VSS VSS nch W=0.8U L=0.24U
M28 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M29 TP8 QN VDD VDD pch W=1.3U L=0.24U
M21 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M9 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M10 TP2 TP21 TP1 VDD pch W=1.3U L=0.24U
M11 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M12 TP2 CLRB TP9 VSS nch W=0.8U L=0.24U
M13 TP9 TP21 VSS VSS nch W=0.8U L=0.24U
M14 TP9 TP0 VSS VSS nch W=0.8U L=0.24U
M7 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M8 TP0 SETB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffss1 SETB DIN SSEL SDIN CLK QN Q
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M8 TP0 SETB VSS VSS nch W=0.8U L=0.24U
M7 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M14 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M15 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M16 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M21 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M23 TP6 CLK TP7 VSS nch W=0.8U L=0.24U
M24 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M29 QN TP7 VDD VDD pch W=3.14U L=0.24U
M30 QN TP7 VSS VSS nch W=2.06U L=0.24U
M17 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M18 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M20 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M25 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M31 Q QN VDD VDD pch W=2.94U L=0.24U
M32 Q QN VSS VSS nch W=1.28U L=0.24U
M22 TP6 TP4 VSS VSS nch W=0.8U L=0.24U
M13 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M28 TP8 QN VSS VSS nch W=0.8U L=0.24U
M11 TP2 TP21 VSS VSS nch W=0.8U L=0.24U
M12 TP2 TP0 VSS VSS nch W=0.8U L=0.24U
M26 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M27 TP8 QN VDD VDD pch W=1.3U L=0.24U
M19 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M9 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M10 TP2 TP21 TP1 VDD pch W=1.3U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sdffss2 SETB DIN SSEL SDIN CLK QN Q
M6 SDIN SSEL TP21 VSS nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M8 TP0 SETB VSS VSS nch W=0.8U L=0.24U
M7 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M14 TP3 CLK VSS VSS nch W=0.8U L=0.24U
M15 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M16 TP2 TP3 TP4 VSS nch W=0.8U L=0.24U
M21 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M23 TP6 CLK TP7 VSS nch W=1.3U L=0.24U
M24 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M29 QN TP7 VDD VDD pch W=6.24U L=0.24U
M30 QN TP7 VSS VSS nch W=3.98U L=0.24U
M17 TP4 CLK TP5 VSS nch W=0.8U L=0.24U
M18 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M20 TP5 TP6 VSS VSS nch W=0.8U L=0.24U
M25 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M31 Q QN VDD VDD pch W=5.92U L=0.24U
M32 Q QN VSS VSS nch W=2.66U L=0.24U
M22 TP6 TP4 VSS VSS nch W=1.26U L=0.24U
M13 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M28 TP8 QN VSS VSS nch W=0.8U L=0.24U
M11 TP2 TP21 VSS VSS nch W=0.8U L=0.24U
M12 TP2 TP0 VSS VSS nch W=0.8U L=0.24U
M26 TP7 TP3 TP8 VSS nch W=0.8U L=0.24U
M27 TP8 QN VDD VDD pch W=1.3U L=0.24U
M19 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL VSS VSS nch W=0.8U L=0.24U
M4 DIN TP20 TP21 VSS nch W=0.8U L=0.24U
M9 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M10 TP2 TP21 TP1 VDD pch W=1.3U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sub1s1 OUTD OUTC0 AIN BIN CIN
M5 N1N303 N1N388 N1N305 VSS nch W=0.8U L=0.24U
M3 N1N301 AIN VDD VDD pch W=1.2U L=0.24U
M4 N1N303 N1N388 N1N301 VDD pch W=1.1U L=0.24U
M7 N1N307 AIN VDD VDD pch W=1.2U L=0.24U
M8 VDD N1N388 N1N307 VDD pch W=1.2U L=0.24U
M9 N1N307 CIN N1N303 VDD pch W=1.1U L=0.24U
M6 N1N305 AIN VSS VSS nch W=0.9U L=0.24U
M10 N1N312 CIN N1N303 VSS nch W=0.8U L=0.24U
M12 VSS N1N388 N1N312 VSS nch W=0.9U L=0.24U
M11 N1N312 AIN VSS VSS nch W=0.9U L=0.24U
M13 N1N337 AIN VDD VDD pch W=1.4U L=0.24U
M17 N1N341 N1N303 N1N337 VDD pch W=1.1U L=0.24U
M14 VDD CIN N1N337 VDD pch W=1.4U L=0.24U
M18 N1N341 N1N303 N1N366 VSS nch W=0.9U L=0.24U
M20 N1N366 CIN VSS VSS nch W=0.9U L=0.24U
M19 N1N366 AIN VSS VSS nch W=0.9U L=0.24U
M21 VSS N1N388 N1N366 VSS nch W=0.9U L=0.24U
M15 VDD N1N388 N1N337 VDD pch W=1.4U L=0.24U
M16 VDD AIN N1N359 VDD pch W=2.1U L=0.24U
M22 N1N359 N1N388 N1N357 VDD pch W=2.1U L=0.24U
M23 N1N357 CIN N1N341 VDD pch W=2.1U L=0.24U
M24 N1N348 CIN N1N341 VSS nch W=1.3U L=0.24U
M25 N1N352 N1N388 N1N348 VSS nch W=1.3U L=0.24U
M26 VSS AIN N1N352 VSS nch W=1.3U L=0.24U
M28 OUTD N1N341 VSS VSS nch W=0.9U L=0.24U
M27 OUTD N1N341 VDD VDD pch W=1.36U L=0.24U
M2 N1N388 BIN VSS VSS nch W=0.6U L=0.24U
M1 N1N388 BIN VDD VDD pch W=1.2U L=0.24U
M30 OUTC0 N1N303 VSS VSS nch W=0.9U L=0.24U
M29 OUTC0 N1N303 VDD VDD pch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sub1s2 OUTD OUTC0 AIN BIN CIN
M5 N1N303 N1N388 N1N305 VSS nch W=1.1U L=0.24U
M3 N1N301 AIN VDD VDD pch W=1.8U L=0.24U
M4 N1N303 N1N388 N1N301 VDD pch W=1.7U L=0.24U
M7 N1N307 AIN VDD VDD pch W=1.8U L=0.24U
M8 VDD N1N388 N1N307 VDD pch W=1.8U L=0.24U
M9 N1N307 CIN N1N303 VDD pch W=1.7U L=0.24U
M6 N1N305 AIN VSS VSS nch W=1.2U L=0.24U
M10 N1N312 CIN N1N303 VSS nch W=1.1U L=0.24U
M12 VSS N1N388 N1N312 VSS nch W=1.2U L=0.24U
M11 N1N312 AIN VSS VSS nch W=1.2U L=0.24U
M13 N1N337 AIN VDD VDD pch W=2.1U L=0.24U
M17 N1N341 N1N303 N1N337 VDD pch W=1.66U L=0.24U
M14 VDD CIN N1N337 VDD pch W=2.1U L=0.24U
M18 N1N341 N1N303 N1N366 VSS nch W=1.16U L=0.24U
M20 N1N366 CIN VSS VSS nch W=1.16U L=0.24U
M19 N1N366 AIN VSS VSS nch W=1.16U L=0.24U
M21 VSS N1N388 N1N366 VSS nch W=1.16U L=0.24U
M15 VDD N1N388 N1N337 VDD pch W=2.1U L=0.24U
M16 VDD AIN N1N359 VDD pch W=3.16U L=0.24U
M22 N1N359 N1N388 N1N357 VDD pch W=3.16U L=0.24U
M23 N1N357 CIN N1N341 VDD pch W=3.16U L=0.24U
M24 N1N348 CIN N1N341 VSS nch W=1.74U L=0.24U
M25 N1N352 N1N388 N1N348 VSS nch W=1.74U L=0.24U
M26 VSS AIN N1N352 VSS nch W=1.74U L=0.24U
M28 OUTD N1N341 VSS VSS nch W=1.44U L=0.24U
M27 OUTD N1N341 VDD VDD pch W=2.48U L=0.24U
M2 N1N388 BIN VSS VSS nch W=0.6U L=0.24U
M1 N1N388 BIN VDD VDD pch W=1.2U L=0.24U
M30 OUTC0 N1N303 VSS VSS nch W=1.46U L=0.24U
M29 OUTC0 N1N303 VDD VDD pch W=2.32U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT sub1s3 OUTD OUTC0 AIN BIN CIN
M5 N1N303 N1N388 N1N305 VSS nch W=1.6U L=0.24U
M3 N1N301 AIN VDD VDD pch W=2.7U L=0.24U
M4 N1N303 N1N388 N1N301 VDD pch W=2.6U L=0.24U
M7 N1N307 AIN VDD VDD pch W=2.7U L=0.24U
M8 VDD N1N388 N1N307 VDD pch W=2.7U L=0.24U
M9 N1N307 CIN N1N303 VDD pch W=2.6U L=0.24U
M6 N1N305 AIN VSS VSS nch W=1.7U L=0.24U
M10 N1N312 CIN N1N303 VSS nch W=1.6U L=0.24U
M12 VSS N1N388 N1N312 VSS nch W=1.7U L=0.24U
M11 N1N312 AIN VSS VSS nch W=1.7U L=0.24U
M13 N1N337 AIN VDD VDD pch W=2.9U L=0.24U
M17 N1N341 N1N303 N1N337 VDD pch W=2.8U L=0.24U
M14 VDD CIN N1N337 VDD pch W=2.9U L=0.24U
M18 N1N341 N1N303 N1N366 VSS nch W=1.52U L=0.24U
M20 N1N366 CIN VSS VSS nch W=1.52U L=0.24U
M19 N1N366 AIN VSS VSS nch W=1.52U L=0.24U
M21 VSS N1N388 N1N366 VSS nch W=1.52U L=0.24U
M15 VDD N1N388 N1N337 VDD pch W=2.9U L=0.24U
M16 VDD AIN N1N359 VDD pch W=4.4U L=0.24U
M22 N1N359 N1N388 N1N357 VDD pch W=4.4U L=0.24U
M23 N1N357 CIN N1N341 VDD pch W=4.3U L=0.24U
M24 N1N348 CIN N1N341 VSS nch W=2.26U L=0.24U
M25 N1N352 N1N388 N1N348 VSS nch W=2.26U L=0.24U
M26 VSS AIN N1N352 VSS nch W=2.26U L=0.24U
M28 OUTD N1N341 VSS VSS nch W=2.9U L=0.24U
M27 OUTD N1N341 VDD VDD pch W=5U L=0.24U
M2 N1N388 BIN VSS VSS nch W=0.7U L=0.24U
M1 N1N388 BIN VDD VDD pch W=1.4U L=0.24U
M30 OUTC0 N1N303 VSS VSS nch W=2.9U L=0.24U
M29 OUTC0 N1N303 VDD VDD pch W=4.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibh1s1 Q E DIN
M2 N1N502 E VSS VSS nch W=0.8U L=0.24U
M1 N1N502 E VDD VDD pch W=1.2U L=0.24U
M5 Q E N1N508 VSS nch W=0.8U L=0.24U
M3 N1N504 DIN VDD VDD pch W=2.3U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=2.3U L=0.24U
M6 N1N508 DIN VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibh1s2 Q E DIN
M2 N1N502 E VSS VSS nch W=0.9U L=0.24U
M1 N1N502 E VDD VDD pch W=1.6U L=0.24U
M5 Q E N1N508 VSS nch W=1U L=0.24U
M3 N1N504 DIN VDD VDD pch W=3U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=3U L=0.24U
M6 N1N508 DIN VSS VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibh1s3 Q E DIN
M2 N1N502 E VSS VSS nch W=1.1U L=0.24U
M1 N1N502 E VDD VDD pch W=2.1U L=0.24U
M5 Q E N1N508 VSS nch W=1.3U L=0.24U
M3 N1N504 DIN VDD VDD pch W=3.9U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=3.9U L=0.24U
M6 N1N508 DIN VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibh1s4 Q E DIN
M2 N1N502 E VSS VSS nch W=2U L=0.24U
M1 N1N502 E VDD VDD pch W=3U L=0.24U
M5 Q E N1N508 VSS nch W=2.1U L=0.24U
M3 N1N504 DIN VDD VDD pch W=6.3U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=6.3U L=0.24U
M6 N1N508 DIN VSS VSS nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibh1s5 Q E DIN
M2 N1N502 E VSS VSS nch W=2.3U L=0.24U
M1 N1N502 E VDD VDD pch W=3.7U L=0.24U
M5 Q E N1N508 VSS nch W=3U L=0.24U
M3 N1N504 DIN VDD VDD pch W=9.32U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=9.32U L=0.24U
M6 N1N508 DIN VSS VSS nch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibh1s6 Q E DIN
M2 N1N502 E VSS VSS nch W=2.9U L=0.24U
M1 N1N502 E VDD VDD pch W=4.8U L=0.24U
M3 N1N504 DIN VDD VDD pch W=11.4U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=11.4U L=0.24U
M5 Q E N1N508 VSS nch W=3.6U L=0.24U
M6 N1N508 DIN VSS VSS nch W=3.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibl1s1 Q EB DIN
M2 N1N510 EB VSS VSS nch W=0.8U L=0.24U
M1 N1N510 EB VDD VDD pch W=1.2U L=0.24U
M3 N1N504 DIN VDD VDD pch W=2.2U L=0.24U
M4 Q EB N1N504 VDD pch W=2.2U L=0.24U
M5 Q N1N510 N1N508 VSS nch W=0.86U L=0.24U
M6 N1N508 DIN VSS VSS nch W=0.86U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibl1s2 Q EB DIN
M2 N1N510 EB VSS VSS nch W=0.9U L=0.24U
M1 N1N510 EB VDD VDD pch W=1.6U L=0.24U
M3 N1N504 DIN VDD VDD pch W=2.8U L=0.24U
M4 Q EB N1N504 VDD pch W=2.8U L=0.24U
M5 Q N1N510 N1N508 VSS nch W=1.16U L=0.24U
M6 N1N508 DIN VSS VSS nch W=1.16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibl1s3 Q EB DIN
M2 N1N510 EB VSS VSS nch W=1.1U L=0.24U
M1 N1N510 EB VDD VDD pch W=2.1U L=0.24U
M3 N1N504 DIN VDD VDD pch W=3.6U L=0.24U
M4 Q EB N1N504 VDD pch W=3.6U L=0.24U
M5 Q N1N510 N1N508 VSS nch W=1.5U L=0.24U
M6 N1N508 DIN VSS VSS nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibl1s4 Q EB DIN
M2 N1N510 EB VSS VSS nch W=1.8U L=0.24U
M1 N1N510 EB VDD VDD pch W=3.5U L=0.24U
M3 N1N504 DIN VDD VDD pch W=5.4U L=0.24U
M4 Q EB N1N504 VDD pch W=5.4U L=0.24U
M5 Q N1N510 N1N508 VSS nch W=2.4U L=0.24U
M6 N1N508 DIN VSS VSS nch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibl1s5 Q EB DIN
M2 N1N510 EB VSS VSS nch W=1.8U L=0.24U
M1 N1N510 EB VDD VDD pch W=3.7U L=0.24U
M3 N1N504 DIN VDD VDD pch W=8.7U L=0.24U
M4 Q EB N1N504 VDD pch W=8.7U L=0.24U
M5 Q N1N510 N1N508 VSS nch W=4.5U L=0.24U
M6 N1N508 DIN VSS VSS nch W=4.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tibl1s6 Q EB DIN
M2 N1N510 EB VSS VSS nch W=2.2U L=0.24U
M1 N1N510 EB VDD VDD pch W=4.4U L=0.24U
M3 N1N504 DIN VDD VDD pch W=11.3U L=0.24U
M4 Q EB N1N504 VDD pch W=11.3U L=0.24U
M5 Q N1N510 N1N508 VSS nch W=6.2U L=0.24U
M6 N1N508 DIN VSS VSS nch W=6.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbh1s1 Q E DIN
M2 N1N517 N1N509 VDD VDD pch W=2.6U L=0.24U
M1 N1N513 E VDD VDD pch W=1.5U L=0.24U
M4 N1N513 E VSS VSS nch W=0.9U L=0.24U
M6 Q E N1N523 VSS nch W=0.94U L=0.24U
M8 N1N523 N1N509 VSS VSS nch W=0.94U L=0.24U
M7 N1N509 DIN VSS VSS nch W=0.8U L=0.24U
M3 Q N1N513 N1N517 VDD pch W=2.6U L=0.24U
M5 N1N509 DIN VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbh1s2 Q E DIN
M2 N1N286 E VSS VSS nch W=0.9U L=0.24U
M1 N1N286 E VDD VDD pch W=1.6U L=0.24U
M4 N1N260 DIN VSS VSS nch W=0.8U L=0.24U
M3 N1N260 DIN VDD VDD pch W=1.6U L=0.24U
M8 N1N267 N1N260 VSS VSS nch W=1.24U L=0.24U
M7 Q E N1N267 VSS nch W=1.24U L=0.24U
M6 Q N1N286 N1N262 VDD pch W=3.6U L=0.24U
M5 N1N262 N1N260 VDD VDD pch W=3.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbh1s3 Q E DIN
M6 N1N565 DIN VDD VDD pch W=1.4U L=0.24U
M1 N1N563 E VDD VDD pch W=1.3U L=0.24U
M3 N1N565 E VDD VDD pch W=1.4U L=0.24U
M9 Q N1N565 VDD VDD pch W=2.42U L=0.24U
M7 N1N567 N1N563 N1N565 VDD pch W=1.3U L=0.24U
M8 N1N567 DIN VSS VSS nch W=0.9U L=0.24U
M10 Q N1N567 VSS VSS nch W=1.46U L=0.24U
M4 N1N565 E N1N567 VSS nch W=0.8U L=0.24U
M2 N1N563 E VSS VSS nch W=0.8U L=0.24U
M5 N1N567 N1N563 VSS VSS nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbh1s4 Q E DIN
M6 N1N565 DIN VDD VDD pch W=2.4U L=0.24U
M1 N1N563 E VDD VDD pch W=1.3U L=0.24U
M3 N1N565 E VDD VDD pch W=2U L=0.24U
M9 Q N1N565 VDD VDD pch W=3.3U L=0.24U
M7 N1N567 N1N563 N1N565 VDD pch W=2.6U L=0.24U
M8 N1N567 DIN VSS VSS nch W=1.2U L=0.24U
M10 Q N1N567 VSS VSS nch W=1.9U L=0.24U
M4 N1N565 E N1N567 VSS nch W=1.4U L=0.24U
M2 N1N563 E VSS VSS nch W=1U L=0.24U
M5 N1N567 N1N563 VSS VSS nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbh1s5 Q E DIN
M6 N1N565 DIN VDD VDD pch W=4U L=0.24U
M1 N1N563 E VDD VDD pch W=3U L=0.24U
M3 N1N565 E VDD VDD pch W=3.1U L=0.24U
M9 Q N1N565 VDD VDD pch W=6.3U L=0.24U
M7 N1N567 N1N563 N1N565 VDD pch W=4.9U L=0.24U
M8 N1N567 DIN VSS VSS nch W=1.4U L=0.24U
M10 Q N1N567 VSS VSS nch W=3.1U L=0.24U
M4 N1N565 E N1N567 VSS nch W=3.1U L=0.24U
M2 N1N563 E VSS VSS nch W=1.8U L=0.24U
M5 N1N567 N1N563 VSS VSS nch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbh1s6 Q E DIN
M6 N1N565 DIN VDD VDD pch W=4.8U L=0.24U
M1 N1N563 E VDD VDD pch W=3.6U L=0.24U
M3 N1N565 E VDD VDD pch W=3.7U L=0.24U
M9 Q N1N565 VDD VDD pch W=7.6U L=0.24U
M7 N1N567 N1N563 N1N565 VDD pch W=5.9U L=0.24U
M8 N1N567 DIN VSS VSS nch W=1.8U L=0.24U
M10 Q N1N567 VSS VSS nch W=3.8U L=0.24U
M4 N1N565 E N1N567 VSS nch W=3.7U L=0.24U
M2 N1N563 E VSS VSS nch W=2.2U L=0.24U
M5 N1N567 N1N563 VSS VSS nch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbl1s1 Q EB DIN
M2 N1N260 DIN VSS VSS nch W=0.9U L=0.24U
M1 N1N260 DIN VDD VDD pch W=1.5U L=0.24U
M4 N1N276 EB VSS VSS nch W=0.8U L=0.24U
M3 N1N276 EB VDD VDD pch W=1.3U L=0.24U
M8 N1N267 N1N260 VSS VSS nch W=0.94U L=0.24U
M7 Q N1N276 N1N267 VSS nch W=0.94U L=0.24U
M6 Q EB N1N262 VDD pch W=2.6U L=0.24U
M5 N1N262 N1N260 VDD VDD pch W=2.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbl1s2 Q EB DIN
M2 N1N260 DIN VSS VSS nch W=0.9U L=0.24U
M1 N1N260 DIN VDD VDD pch W=1.6U L=0.24U
M4 N1N276 EB VSS VSS nch W=0.9U L=0.24U
M3 N1N276 EB VDD VDD pch W=1.8U L=0.24U
M8 N1N267 N1N260 VSS VSS nch W=1.26U L=0.24U
M7 Q N1N276 N1N267 VSS nch W=1.26U L=0.24U
M6 Q EB N1N262 VDD pch W=3.5U L=0.24U
M5 N1N262 N1N260 VDD VDD pch W=3.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbl1s3 Q EB DIN
M4 N1N259 DIN VSS VSS nch W=1.9U L=0.24U
M2 N1N257 DIN VDD VDD pch W=1.5U L=0.24U
M3 N1N259 EB N1N257 VDD pch W=1.6U L=0.24U
M5 N1N257 N1N285 VDD VDD pch W=1U L=0.24U
M6 N1N257 N1N285 N1N259 VSS nch W=1.5U L=0.24U
M7 N1N259 EB VSS VSS nch W=1U L=0.24U
M9 Q N1N259 VSS VSS nch W=1.46U L=0.24U
M8 Q N1N257 VDD VDD pch W=2.42U L=0.24U
M1 N1N285 EB VDD VDD pch W=1.3U L=0.24U
M10 N1N285 EB VSS VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbl1s4 Q EB DIN
M4 N1N259 DIN VSS VSS nch W=2.5U L=0.24U
M2 N1N257 DIN VDD VDD pch W=2.8U L=0.24U
M3 N1N259 EB N1N257 VDD pch W=2.8U L=0.24U
M5 N1N257 N1N285 VDD VDD pch W=1.7U L=0.24U
M6 N1N257 N1N285 N1N259 VSS nch W=1.8U L=0.24U
M7 N1N259 EB VSS VSS nch W=1.6U L=0.24U
M9 Q N1N259 VSS VSS nch W=1.92U L=0.24U
M8 Q N1N257 VDD VDD pch W=4U L=0.24U
M1 N1N285 EB VDD VDD pch W=1.7U L=0.24U
M10 N1N285 EB VSS VSS nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbl1s5 Q EB DIN
M4 N1N259 DIN VSS VSS nch W=3.1U L=0.24U
M2 N1N257 DIN VDD VDD pch W=3.5U L=0.24U
M3 N1N259 EB N1N257 VDD pch W=3.8U L=0.24U
M5 N1N257 N1N285 VDD VDD pch W=2.1U L=0.24U
M6 N1N257 N1N285 N1N259 VSS nch W=2.2U L=0.24U
M7 N1N259 EB VSS VSS nch W=1.6U L=0.24U
M9 Q N1N259 VSS VSS nch W=3.1U L=0.24U
M8 Q N1N257 VDD VDD pch W=7U L=0.24U
M1 N1N285 EB VDD VDD pch W=2.2U L=0.24U
M10 N1N285 EB VSS VSS nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT tnbl1s6 Q EB DIN
M4 N1N259 DIN VSS VSS nch W=3.7U L=0.24U
M2 N1N257 DIN VDD VDD pch W=4.2U L=0.24U
M3 N1N259 EB N1N257 VDD pch W=4.6U L=0.24U
M5 N1N257 N1N285 VDD VDD pch W=2.5U L=0.24U
M6 N1N257 N1N285 N1N259 VSS nch W=2.6U L=0.24U
M7 N1N259 EB VSS VSS nch W=1.9U L=0.24U
M9 Q N1N259 VSS VSS nch W=3.7U L=0.24U
M8 Q N1N257 VDD VDD pch W=8.6U L=0.24U
M1 N1N285 EB VDD VDD pch W=2.6U L=0.24U
M10 N1N285 EB VSS VSS nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xnr2s1 Q DIN1 DIN2
M9 Q N1N89 VDD VDD pch W=3.1U L=0.24U 
M10 Q N1N89 VSS VSS nch W=1.1U L=0.24U 
M4 N1N123 DIN1 VSS VSS nch W=0.6U L=0.24U 
M3 N1N123 DIN1 VDD VDD pch W=1.5U L=0.24U 
M2 N1N83 DIN2 VSS VSS nch W=0.6U L=0.24U 
M1 N1N83 DIN2 VDD VDD pch W=1.3U L=0.24U 
M5 N1N89 DIN1 DIN2 VDD pch W=1.4U L=0.24U 
M6 DIN2 N1N123 N1N89 VSS nch W=0.6U L=0.24U 
M8 N1N83 DIN1 N1N89 VSS nch W=0.6U L=0.24U 
M7 N1N89 N1N123 N1N83 VDD pch W=1.4U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xnr2s2 Q DIN1 DIN2
M10 Q N1N89 VSS VSS nch W=2.2U L=0.24U 
M4 N1N83 DIN1 VSS VSS nch W=1.2U L=0.24U 
M3 N1N83 DIN1 VDD VDD pch W=3U L=0.24U 
M2 N1N121 DIN2 VSS VSS nch W=1.5U L=0.24U 
M1 N1N121 DIN2 VDD VDD pch W=2.8U L=0.24U 
M5 N1N89 DIN1 DIN2 VDD pch W=2U L=0.24U 
M6 DIN2 N1N83 N1N89 VSS nch W=0.8U L=0.24U 
M8 N1N121 DIN1 N1N89 VSS nch W=0.8U L=0.24U 
M7 N1N89 N1N83 N1N121 VDD pch W=2U L=0.24U 
M9 Q N1N89 VDD VDD pch W=5.5U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xnr2s3 Q DIN1 DIN2
M10 Q N1N89 VSS VSS nch W=3.8U L=0.24U 
M4 N1N83 DIN1 VSS VSS nch W=2.4U L=0.24U 
M3 N1N83 DIN1 VDD VDD pch W=5.8U L=0.24U 
M2 N1N121 DIN2 VSS VSS nch W=2.9U L=0.24U 
M1 N1N121 DIN2 VDD VDD pch W=5.2U L=0.24U 
M5 N1N89 DIN1 DIN2 VDD pch W=3U L=0.24U 
M6 DIN2 N1N83 N1N89 VSS nch W=1.2U L=0.24U 
M8 N1N121 DIN1 N1N89 VSS nch W=1.2U L=0.24U 
M7 N1N89 N1N83 N1N121 VDD pch W=3U L=0.24U 
M9 Q N1N89 VDD VDD pch W=9.5U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xnr3s1 Q DIN1 DIN2 DIN3
M20 Q N1N299 VSS VSS nch W=2.9U L=0.24U 
M19 Q N1N299 VDD VDD pch W=3.8U L=0.24U 
M15 N1N299 N1N328 DIN2 VDD pch W=1.5U L=0.24U 
M16 DIN2 N1N321 N1N299 VSS nch W=0.6U L=0.24U 
M2 N1N309 DIN1 VSS VSS nch W=1.1U L=0.24U 
M1 N1N309 DIN1 VDD VDD pch W=2.6U L=0.24U 
M4 N1N313 DIN2 VSS VSS nch W=0.6U L=0.24U 
M3 N1N313 DIN2 VDD VDD pch W=1.8U L=0.24U 
M6 N1N317 DIN3 VSS VSS nch W=1.2U L=0.24U 
M5 N1N317 DIN3 VDD VDD pch W=2.4U L=0.24U 
M8 N1N317 N1N309 N1N321 VSS nch W=0.7U L=0.24U 
M7 N1N321 DIN1 N1N317 VDD pch W=1.7U L=0.24U 
M10 DIN3 DIN1 N1N321 VSS nch W=0.7U L=0.24U 
M9 N1N321 N1N309 DIN3 VDD pch W=1.7U L=0.24U 
M11 N1N328 DIN1 DIN3 VDD pch W=1.7U L=0.24U 
M12 DIN3 N1N309 N1N328 VSS nch W=0.7U L=0.24U 
M13 N1N328 N1N309 N1N317 VDD pch W=1.7U L=0.24U 
M14 N1N317 DIN1 N1N328 VSS nch W=0.7U L=0.24U 
M18 N1N313 N1N328 N1N299 VSS nch W=0.6U L=0.24U 
M17 N1N299 N1N321 N1N313 VDD pch W=1.5U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xnr3s2 Q DIN1 DIN2 DIN3
M20 Q N1N299 VSS VSS nch W=4.4U L=0.24U 
M19 Q N1N299 VDD VDD pch W=5.7U L=0.24U 
M15 N1N299 N1N328 DIN2 VDD pch W=2.1U L=0.24U 
M16 DIN2 N1N321 N1N299 VSS nch W=0.8U L=0.24U 
M2 N1N309 DIN1 VSS VSS nch W=1.7U L=0.24U 
M1 N1N309 DIN1 VDD VDD pch W=3.9U L=0.24U 
M4 N1N313 DIN2 VSS VSS nch W=1U L=0.24U 
M3 N1N313 DIN2 VDD VDD pch W=2.6U L=0.24U 
M6 N1N317 DIN3 VSS VSS nch W=1.8U L=0.24U 
M5 N1N317 DIN3 VDD VDD pch W=3.6U L=0.24U 
M8 N1N317 N1N309 N1N321 VSS nch W=1U L=0.24U 
M7 N1N321 DIN1 N1N317 VDD pch W=2.4U L=0.24U 
M10 DIN3 DIN1 N1N321 VSS nch W=1U L=0.24U 
M9 N1N321 N1N309 DIN3 VDD pch W=2.4U L=0.24U 
M11 N1N328 DIN1 DIN3 VDD pch W=2.4U L=0.24U 
M12 DIN3 N1N309 N1N328 VSS nch W=1U L=0.24U 
M13 N1N328 N1N309 N1N317 VDD pch W=2.4U L=0.24U 
M14 N1N317 DIN1 N1N328 VSS nch W=1U L=0.24U 
M18 N1N313 N1N328 N1N299 VSS nch W=0.8U L=0.24U 
M17 N1N299 N1N321 N1N313 VDD pch W=2.1U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xnr3s3 Q DIN1 DIN2 DIN3
M20 Q N1N299 VSS VSS nch W=7.1U L=0.24U 
M19 Q N1N299 VDD VDD pch W=9.5U L=0.24U 
M15 N1N299 N1N328 DIN2 VDD pch W=3.2U L=0.24U 
M16 DIN2 N1N321 N1N299 VSS nch W=1.2U L=0.24U 
M2 N1N309 DIN1 VSS VSS nch W=3.1U L=0.24U 
M1 N1N309 DIN1 VDD VDD pch W=7U L=0.24U 
M4 N1N313 DIN2 VSS VSS nch W=1.8U L=0.24U 
M3 N1N313 DIN2 VDD VDD pch W=4.4U L=0.24U 
M6 N1N317 DIN3 VSS VSS nch W=3.2U L=0.24U 
M5 N1N317 DIN3 VDD VDD pch W=6.5U L=0.24U 
M8 N1N317 N1N309 N1N321 VSS nch W=1.5U L=0.24U 
M7 N1N321 DIN1 N1N317 VDD pch W=3.6U L=0.24U 
M10 DIN3 DIN1 N1N321 VSS nch W=1.5U L=0.24U 
M9 N1N321 N1N309 DIN3 VDD pch W=3.6U L=0.24U 
M11 N1N328 DIN1 DIN3 VDD pch W=3.6U L=0.24U 
M12 DIN3 N1N309 N1N328 VSS nch W=1.5U L=0.24U 
M13 N1N328 N1N309 N1N317 VDD pch W=3.6U L=0.24U 
M14 N1N317 DIN1 N1N328 VSS nch W=1.5U L=0.24U 
M18 N1N313 N1N328 N1N299 VSS nch W=1.2U L=0.24U 
M17 N1N299 N1N321 N1N313 VDD pch W=3.2U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xor2s1 Q DIN1 DIN2
M2       N1N83 DIN1 VSS    VSS nch W=0.6U L=0.24U
M1       N1N83 DIN1 VDD  VDD pch W=1.3U L=0.24U
M4       N1N85 DIN2 VSS    VSS nch W=0.6U L=0.24U
M3       N1N85 DIN2 VDD  VDD pch W=1.5U L=0.24U
M5       N1N91 DIN2 N1N83  VDD pch W=1.4U L=0.24U
M6       N1N83 N1N85 N1N91  VSS nch W=0.6U L=0.24U
M8       DIN1 DIN2 N1N91  VSS nch W=0.6U L=0.24U
M7       N1N91 N1N85 DIN1  VDD pch W=1.4U L=0.24U
M10      Q N1N91 VSS    VSS nch W=1.9U L=0.24U
M9       Q N1N91 VDD  VDD pch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xor2s2 Q DIN1 DIN2
M2       N1N83 DIN1 VSS    VSS nch W=1.2U L=0.24U
M1       N1N83 DIN1 VDD  VDD pch W=2.6U L=0.24U
M4       N1N85 DIN2 VSS    VSS nch W=1.2U L=0.24U
M3       N1N85 DIN2 VDD  VDD pch W=3.0U L=0.24U
M5       N1N91 DIN2 N1N83  VDD pch W=2.0U L=0.24U
M6       N1N83 N1N85 N1N91  VSS nch W=0.8U L=0.24U
M8       DIN1 DIN2 N1N91  VSS nch W=0.8U L=0.24U
M7       N1N91 N1N85 DIN1  VDD pch W=2.0U L=0.24U
M10      Q N1N91 VSS    VSS nch W=3.7U L=0.24U
M9       Q N1N91 VDD  VDD pch W=5.0U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xor2s3 Q DIN1 DIN2
M2       N1N83 DIN1 VSS    VSS nch W=2.4U L=0.24U
M1       N1N83 DIN1 VDD  VDD pch W=5.2U L=0.24U
M4       N1N85 DIN2 VSS    VSS nch W=2.4U L=0.24U
M3       N1N85 DIN2 VDD  VDD pch W=5.8U L=0.24U
M5       N1N91 DIN2 N1N83  VDD pch W=3.0U L=0.24U
M6       N1N83 N1N85 N1N91  VSS nch W=1.2U L=0.24U
M8       DIN1 DIN2 N1N91  VSS nch W=1.2U L=0.24U
M7       N1N91 N1N85 DIN1  VDD pch W=3.0U L=0.24U
M10      Q N1N91 VSS    VSS nch W=6.7U L=0.24U
M9       Q N1N91 VDD  VDD pch W=9.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xor3s1 Q DIN1 DIN2 DIN3
M20      Q N1N307 VSS    VSS nch W=2.9U L=0.24U
M19      Q N1N307 VDD  VDD pch W=3.8U L=0.24U
M15      N1N307 DIN2 N1N311  VDD pch W=1.5U L=0.24U
M16      N1N311 N1N321 N1N307  VSS nch W=0.6U L=0.24U
M2       N1N360 DIN1 VSS    VSS nch W=1.1U L=0.24U
M1       N1N360 DIN1 VDD  VDD pch W=2.6U L=0.24U
M4       N1N321 DIN2 VSS    VSS nch W=0.7U L=0.24U
M3       N1N321 DIN2 VDD  VDD pch W=1.4U L=0.24U
M6       N1N325 DIN3 VSS    VSS nch W=1.2U L=0.24U
M5       N1N325 DIN3 VDD  VDD pch W=2.4U L=0.24U
M7       N1N311 DIN1 N1N325  VDD pch W=1.7U L=0.24U
M8       N1N325 N1N360 N1N311  VSS nch W=0.7U L=0.24U
M10      DIN3 DIN1 N1N311  VSS nch W=0.7U L=0.24U
M9       N1N311 N1N360 DIN3  VDD pch W=1.7U L=0.24U
M12      DIN3 N1N360 N1N338  VSS nch W=0.7U L=0.24U
M11      N1N338 DIN1 DIN3  VDD pch W=1.7U L=0.24U
M13      N1N338 N1N360 N1N325  VDD pch W=1.7U L=0.24U
M14      N1N325 DIN1 N1N338  VSS nch W=0.7U L=0.24U
M17      N1N307 N1N321 N1N338  VDD pch W=1.5U L=0.24U
M18      N1N338 DIN2 N1N307  VSS nch W=0.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xor3s2 Q DIN1 DIN2 DIN3
M20      Q N1N307 VSS    VSS nch W=4.4U L=0.24U
M19      Q N1N307 VDD  VDD pch W=5.7U L=0.24U
M15      N1N307 DIN2 N1N311  VDD pch W=2.1U L=0.24U
M16      N1N311 N1N321 N1N307  VSS nch W=0.8U L=0.24U
M2       N1N360 DIN1 VSS    VSS nch W=1.7U L=0.24U
M1       N1N360 DIN1 VDD  VDD pch W=3.9U L=0.24U
M4       N1N321 DIN2 VSS    VSS nch W=1.1U L=0.24U
M3       N1N321 DIN2 VDD  VDD pch W=2.1U L=0.24U
M6       N1N325 DIN3 VSS    VSS nch W=1.8U L=0.24U
M5       N1N325 DIN3 VDD  VDD pch W=3.6U L=0.24U
M7       N1N311 DIN1 N1N325  VDD pch W=2.4U L=0.24U
M8       N1N325 N1N360 N1N311  VSS nch W=1.0U L=0.24U
M10      DIN3 DIN1 N1N311  VSS nch W=1.0U L=0.24U
M9       N1N311 N1N360 DIN3  VDD pch W=2.4U L=0.24U
M12      DIN3 N1N360 N1N338  VSS nch W=1.0U L=0.24U
M11      N1N338 DIN1 DIN3  VDD pch W=2.4U L=0.24U
M13      N1N338 N1N360 N1N325  VDD pch W=2.4U L=0.24U
M14      N1N325 DIN1 N1N338  VSS nch W=1.0U L=0.24U
M17      N1N307 N1N321 N1N338  VDD pch W=2.1U L=0.24U
M18      N1N338 DIN2 N1N307  VSS nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT xor3s3 Q DIN1 DIN2 DIN3
M20      Q N1N307 VSS    VSS nch W=7.1U L=0.24U
M19      Q N1N307 VDD  VDD pch W=9.54U L=0.24U
M15      N1N307 DIN2 N1N311  VDD pch W=3.2U L=0.24U
M16      N1N311 N1N321 N1N307  VSS nch W=1.2U L=0.24U
M2       N1N360 DIN1 VSS    VSS nch W=3.1U L=0.24U
M1       N1N360 DIN1 VDD  VDD pch W=7.0U L=0.24U
M4       N1N321 DIN2 VSS    VSS nch W=2.0U L=0.24U
M3       N1N321 DIN2 VDD  VDD pch W=3.8U L=0.24U
M6       N1N325 DIN3 VSS    VSS nch W=3.2U L=0.24U
M5       N1N325 DIN3 VDD  VDD pch W=6.5U L=0.24U
M7       N1N311 DIN1 N1N325  VDD pch W=3.6U L=0.24U
M8       N1N325 N1N360 N1N311  VSS nch W=1.5U L=0.24U
M10      DIN3 DIN1 N1N311  VSS nch W=1.5U L=0.24U
M9       N1N311 N1N360 DIN3  VDD pch W=3.6U L=0.24U
M12      DIN3 N1N360 N1N338  VSS nch W=1.5U L=0.24U
M11      N1N338 DIN1 DIN3  VDD pch W=3.6U L=0.24U
M13      N1N338 N1N360 N1N325  VDD pch W=3.6U L=0.24U
M14      N1N325 DIN1 N1N338  VSS nch W=1.5U L=0.24U
M17      N1N307 N1N321 N1N338  VDD pch W=3.2U L=0.24U
M18      N1N338 DIN2 N1N307  VSS nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT avdd PAD AVDD
C1I4110 PAD N1I41TP0 235FF
C1I4111 N1I41TP2 PAD 235FF
M1 AVDD N1N17 AVSS AVSS nch W=300U L=0.34U
M1I410 N1I41TP7 N1I41TP0 NVDD NVDD pch W=38U L=0.34U
M1I411 N1I41TP0 N1I41TP1 NVDD NVDD pch W=6U L=6U
M1I412 N1I41TP2 N1I41TP3 NVSS NVSS nch W=6U L=6U
M1I413 N1I41TP4 N1I41TP2 N1I41TP5 NVSS nch W=38U L=0.34U
R1 N1N17 AVSS 400
R1I414 N1I41TP7 EVSS 123
R1I415 NVDD N1I41TP3 198
R1I416 EVDD N1I41TP4 177
R1I417 N1I41TP1 NVSS 198
R1I418 N1I41TP5 NVSS 0.21
R1I419 N1I41TP5 NVSS 0.21
R2 AVDD PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT avss PAD AVSS
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 AVSS N1N48 AVDD AVDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 AVDD N1N48 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 AVSS PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cainr25s4 PAD Q
C1I35710 PAD N1I357TP0 235FF
C1I35711 N1I357TP2 PAD 235FF
M1I3570 N1I357TP7 N1I357TP0 NVDD NVDD pch W=38U L=0.34U
M1I3571 N1I357TP0 N1I357TP1 NVDD NVDD pch W=6U L=6U
M1I3572 N1I357TP2 N1I357TP3 NVSS NVSS nch W=6U L=6U
M1I3573 N1I357TP4 N1I357TP2 N1I357TP5 NVSS nch W=38U L=0.34U
R1 PAD Q 200
R1I3574 N1I357TP7 EVSS 123
R1I3575 NVDD N1I357TP3 198
R1I3576 EVDD N1I357TP4 177
R1I3577 N1I357TP1 NVSS 198
R1I3578 N1I357TP5 NVSS 0.21
R1I3579 N1I357TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT caon25s4 PAD DIN
C1I36910 PAD N1I369TP0 235FF
C1I36911 N1I369TP2 PAD 235FF
M1I3690 N1I369TP7 N1I369TP0 NVDD NVDD pch W=38U L=0.34U
M1I3691 N1I369TP0 N1I369TP1 NVDD NVDD pch W=6U L=6U
M1I3692 N1I369TP2 N1I369TP3 NVSS NVSS nch W=6U L=6U
M1I3693 N1I369TP4 N1I369TP2 N1I369TP5 NVSS nch W=38U L=0.34U
R1 PAD DIN 0.30
R1I3694 N1I369TP7 EVSS 123
R1I3695 NVDD N1I369TP3 198
R1I3696 EVDD N1I369TP4 177
R1I3697 N1I369TP1 NVSS 198
R1I3698 N1I369TP5 NVSS 0.21
R1I3699 N1I369TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cdavdd AVDD PAD VDD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 VDD N1N17 VSS VSS nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N17 VSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 VDD PAD 0.002
R3 AVDD VDD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cdavss AVSS PAD VSS
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 VSS N1N48 VDD VDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 VDD N1N48 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 VSS PAD 0.002
R3 AVSS VSS 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cdvdd PAD VDD N1
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 VDD N1N17 VSS VSS nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N17 VSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 VDD PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cdvss PAD VSS N1
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 VSS N1N48 VDD VDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 VDD N1N48 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 VSS PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cii25s1 PAD Q
C1I38610 PAD N1I386TP0 235FF
C1I38611 N1I386TP2 PAD 235FF
M1 Q TP2 VDD VDD pch W=3.8U L=0.24U
M1I3860 N1I386TP7 N1I386TP0 NVDD NVDD pch W=38U L=0.34U
M1I3861 N1I386TP0 N1I386TP1 NVDD NVDD pch W=6U L=6U
M1I3862 N1I386TP2 N1I386TP3 NVSS NVSS nch W=6U L=6U
M1I3863 N1I386TP4 N1I386TP2 N1I386TP5 NVSS nch W=38U L=0.34U
M2 Q TP2 VSS VSS nch W=1.36U L=0.24U
M6 TP2 VDD VDD VDD pch W=100U L=0.48U
M7 TP2 VSS VSS VSS nch W=100U L=0.48U
R1 TP2 PAD 300
R1I3864 N1I386TP7 EVSS 123
R1I3865 NVDD N1I386TP3 198
R1I3866 EVDD N1I386TP4 177
R1I3867 N1I386TP1 NVSS 198
R1I3868 N1I386TP5 NVSS 0.21
R1I3869 N1I386TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cii25s4 PAD Q
C1I39610 PAD N1I396TP0 235FF
C1I39611 N1I396TP2 PAD 235FF
M1 Q TP2 VDD VDD pch W=30U L=0.24U
M1I3960 N1I396TP7 N1I396TP0 NVDD NVDD pch W=38U L=0.34U
M1I3961 N1I396TP0 N1I396TP1 NVDD NVDD pch W=6U L=6U
M1I3962 N1I396TP2 N1I396TP3 NVSS NVSS nch W=6U L=6U
M1I3963 N1I396TP4 N1I396TP2 N1I396TP5 NVSS nch W=38U L=0.34U
M2 Q TP2 VSS VSS nch W=10.12U L=0.24U
M6 TP2 VDD VDD VDD pch W=100U L=0.48U
M7 TP2 VSS VSS VSS nch W=100U L=0.48U
R1 TP2 PAD 300
R1I3964 N1I396TP7 EVSS 123
R1I3965 NVDD N1I396TP3 198
R1I3966 EVDD N1I396TP4 177
R1I3967 N1I396TP1 NVSS 198
R1I3968 N1I396TP5 NVSS 0.21
R1I3969 N1I396TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ciis25s1 PAD Q
C1I50810 PAD N1I508TP0 235FF
C1I50811 N1I508TP2 PAD 235FF
M1 TP0 TP5 VDD VDD pch W=2.74U L=0.24U
M1I5080 N1I508TP7 N1I508TP0 NVDD NVDD pch W=38U L=0.34U
M1I5081 N1I508TP0 N1I508TP1 NVDD NVDD pch W=6U L=6U
M1I5082 N1I508TP2 N1I508TP3 NVSS NVSS nch W=6U L=6U
M1I5083 N1I508TP4 N1I508TP2 N1I508TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP5 TP0 VDD pch W=2.74U L=0.24U
M3 TP1 TP5 TP2 VSS nch W=24U L=0.24U
M4 TP2 TP5 VSS VSS nch W=24U L=0.24U
M5 VSS TP1 TP0 VDD pch W=7.8U L=0.24U
M6 TP2 TP1 VDD VSS nch W=0.4U L=0.24U
M7 TP3 TP1 VDD VDD pch W=1U L=0.24U
M8 TP3 TP1 VSS VSS nch W=8.2U L=0.24U
M9 Q TP3 VDD VDD pch W=17.5U L=0.24U
M10 Q TP3 VSS VSS nch W=1U L=0.24U
M13 TP5 VDD VDD VDD pch W=100U L=0.48U
M14 TP5 VSS VSS VSS nch W=100U L=0.48U
R1 PAD TP5 300
R1I5084 N1I508TP7 EVSS 123
R1I5085 NVDD N1I508TP3 198
R1I5086 EVDD N1I508TP4 177
R1I5087 N1I508TP1 NVSS 198
R1I5088 N1I508TP5 NVSS 0.21
R1I5089 N1I508TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ciis25s4 PAD Q
C1I49710 PAD N1I497TP0 235FF
C1I49711 N1I497TP2 PAD 235FF
M1 TP0 TP5 VDD VDD pch W=2.74U L=0.24U
M1I4970 N1I497TP7 N1I497TP0 NVDD NVDD pch W=38U L=0.34U
M1I4971 N1I497TP0 N1I497TP1 NVDD NVDD pch W=6U L=6U
M1I4972 N1I497TP2 N1I497TP3 NVSS NVSS nch W=6U L=6U
M1I4973 N1I497TP4 N1I497TP2 N1I497TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP5 TP0 VDD pch W=2.74U L=0.24U
M3 TP1 TP5 TP2 VSS nch W=42U L=0.24U
M4 TP2 TP5 VSS VSS nch W=42U L=0.24U
M5 VSS TP1 TP0 VDD pch W=4.8U L=0.24U
M6 TP2 TP1 VDD VSS nch W=0.4U L=0.24U
M7 TP3 TP1 VDD VDD pch W=1U L=0.24U
M8 TP3 TP1 VSS VSS nch W=8.5U L=0.24U
M9 Q TP3 VDD VDD pch W=15.2U L=0.24U
M10 Q TP3 VSS VSS nch W=1.1U L=0.24U
M13 TP5 VDD VDD VDD pch W=100U L=0.48U
M14 TP5 VSS VSS VSS nch W=100U L=0.48U
R1 PAD TP5 300
R1I4974 N1I497TP7 EVSS 123
R1I4975 NVDD N1I497TP3 198
R1I4976 EVDD N1I497TP4 177
R1I4977 N1I497TP1 NVSS 198
R1I4978 N1I497TP5 NVSS 0.21
R1I4979 N1I497TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cin25s1 PAD Q
C1I38610 PAD N1I386TP0 235FF
C1I38611 N1I386TP2 PAD 235FF
M1 TP1 TP2 VDD VDD pch W=3.8U L=0.24U
M1I3860 N1I386TP7 N1I386TP0 NVDD NVDD pch W=38U L=0.34U
M1I3861 N1I386TP0 N1I386TP1 NVDD NVDD pch W=6U L=6U
M1I3862 N1I386TP2 N1I386TP3 NVSS NVSS nch W=6U L=6U
M1I3863 N1I386TP4 N1I386TP2 N1I386TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP2 VSS VSS nch W=1.36U L=0.24U
M3 Q TP1 VDD VDD pch W=5.6U L=0.24U
M4 Q TP1 VSS VSS nch W=2.6U L=0.24U
M6 TP2 VDD VDD VDD pch W=100U L=0.48U
M7 TP2 VSS VSS VSS nch W=100U L=0.48U
R1 TP2 PAD 300
R1I3864 N1I386TP7 EVSS 123
R1I3865 NVDD N1I386TP3 198
R1I3866 EVDD N1I386TP4 177
R1I3867 N1I386TP1 NVSS 198
R1I3868 N1I386TP5 NVSS 0.21
R1I3869 N1I386TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cin25s4 PAD Q
C1I39610 PAD N1I396TP0 235FF
C1I39611 N1I396TP2 PAD 235FF
M1 TP1 TP2 VDD VDD pch W=30U L=0.24U
M1I3960 N1I396TP7 N1I396TP0 NVDD NVDD pch W=38U L=0.34U
M1I3961 N1I396TP0 N1I396TP1 NVDD NVDD pch W=6U L=6U
M1I3962 N1I396TP2 N1I396TP3 NVSS NVSS nch W=6U L=6U
M1I3963 N1I396TP4 N1I396TP2 N1I396TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP2 VSS VSS nch W=10.12U L=0.24U
M3 Q TP1 VDD VDD pch W=35.52U L=0.24U
M4 Q TP1 VSS VSS nch W=15.92U L=0.24U
M6 TP2 VDD VDD VDD pch W=100U L=0.48U
M7 TP2 VSS VSS VSS nch W=100U L=0.48U
R1 TP2 PAD 300
R1I3964 N1I396TP7 EVSS 123
R1I3965 NVDD N1I396TP3 198
R1I3966 EVDD N1I396TP4 177
R1I3967 N1I396TP1 NVSS 198
R1I3968 N1I396TP5 NVSS 0.21
R1I3969 N1I396TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cins25s1 PAD Q
C1I50810 PAD N1I508TP0 235FF
C1I50811 N1I508TP2 PAD 235FF
M1 TP0 TP5 VDD VDD pch W=2.74U L=0.24U
M1I5080 N1I508TP7 N1I508TP0 NVDD NVDD pch W=38U L=0.34U
M1I5081 N1I508TP0 N1I508TP1 NVDD NVDD pch W=6U L=6U
M1I5082 N1I508TP2 N1I508TP3 NVSS NVSS nch W=6U L=6U
M1I5083 N1I508TP4 N1I508TP2 N1I508TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP5 TP0 VDD pch W=2.74U L=0.24U
M3 TP1 TP5 TP2 VSS nch W=24U L=0.24U
M4 TP2 TP5 VSS VSS nch W=24U L=0.24U
M5 VSS TP1 TP0 VDD pch W=7.8U L=0.24U
M6 TP2 TP1 VDD VSS nch W=0.4U L=0.24U
M7 TP3 TP1 VDD VDD pch W=1U L=0.24U
M8 TP3 TP1 VSS VSS nch W=8.2U L=0.24U
M9 TP4 TP3 VDD VDD pch W=17.5U L=0.24U
M10 TP4 TP3 VSS VSS nch W=1U L=0.24U
M11 Q TP4 VDD VDD pch W=8.2U L=0.24U
M12 Q TP4 VSS VSS nch W=4.1U L=0.24U
M13 TP5 VDD VDD VDD pch W=100U L=0.48U
M14 TP5 VSS VSS VSS nch W=100U L=0.48U
R1 PAD TP5 300
R1I5084 N1I508TP7 EVSS 123
R1I5085 NVDD N1I508TP3 198
R1I5086 EVDD N1I508TP4 177
R1I5087 N1I508TP1 NVSS 198
R1I5088 N1I508TP5 NVSS 0.21
R1I5089 N1I508TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cins25s4 PAD Q
C1I49510 PAD N1I495TP0 235FF
C1I49511 N1I495TP2 PAD 235FF
M1 TP0 TP5 VDD VDD pch W=2.74U L=0.24U
M1I4950 N1I495TP7 N1I495TP0 NVDD NVDD pch W=38U L=0.34U
M1I4951 N1I495TP0 N1I495TP1 NVDD NVDD pch W=6U L=6U
M1I4952 N1I495TP2 N1I495TP3 NVSS NVSS nch W=6U L=6U
M1I4953 N1I495TP4 N1I495TP2 N1I495TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP5 TP0 VDD pch W=2.74U L=0.24U
M3 TP1 TP5 TP2 VSS nch W=42U L=0.24U
M4 TP2 TP5 VSS VSS nch W=42U L=0.24U
M5 VSS TP1 TP0 VDD pch W=4.8U L=0.24U
M6 TP2 TP1 VDD VSS nch W=0.4U L=0.24U
M7 TP3 TP1 VDD VDD pch W=1U L=0.24U
M8 TP3 TP1 VSS VSS nch W=8.5U L=0.24U
M9 TP4 TP3 VDD VDD pch W=15.2U L=0.24U
M10 TP4 TP3 VSS VSS nch W=1.1U L=0.24U
M11 Q TP4 VDD VDD pch W=30.1U L=0.24U
M12 Q TP4 VSS VSS nch W=18.5U L=0.24U
M13 TP5 VDD VDD VDD pch W=100U L=0.48U
M14 TP5 VSS VSS VSS nch W=100U L=0.48U
R1 PAD TP5 300
R1I4954 N1I495TP7 EVSS 123
R1I4955 NVDD N1I495TP3 198
R1I4956 EVDD N1I495TP4 177
R1I4957 N1I495TP1 NVSS 198
R1I4958 N1I495TP5 NVSS 0.21
R1I4959 N1I495TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cioit25s1 DIN E PAD Q
C1I35310 PAD N1I353TP0 235FF
C1I35311 N1I353TP2 PAD 235FF
M1I3530 N1I353TP7 N1I353TP0 NVDD NVDD pch W=38U L=0.34U
M1I3531 N1I353TP0 N1I353TP1 NVDD NVDD pch W=6U L=6U
M1I3532 N1I353TP2 N1I353TP3 NVSS NVSS nch W=6U L=6U
M1I3533 N1I353TP4 N1I353TP2 N1I353TP5 NVSS nch W=38U L=0.34U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E VSS VSS nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=13U L=0.24U
M6 TP2 E TP3 VSS nch W=10U L=0.24U
M7 TP3 TP1 VSS VSS nch W=7U L=0.24U
M8 VDD TP20 TP2 VDD pch W=13U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 VSS TP20 TP3 VSS nch W=7U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=15.5U L=0.34U
M14 TP14 TP3 NVSS VSS nch W=5U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=15.5U L=0.34U
M18 TP15 TP3 NVSS VSS nch W=5U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=15.5U L=0.34U
M22 TP16 TP3 NVSS VSS nch W=5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=15.5U L=0.34U
M26 TP17 TP3 NVSS VSS nch W=5U L=0.34U
M27 PAD NVSS NVSS VSS nch W=34U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 VSS TP4 Q VSS nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 VSS TP13 TP4 VSS nch W=4.1U L=0.24U
M33 TP20 DIN VDD VDD pch W=5.4U L=0.24U
M34 TP20 DIN VSS VSS nch W=7U L=0.24U
R1I3534 N1I353TP7 EVSS 123
R1I3535 NVDD N1I353TP3 198
R1I3536 EVDD N1I353TP4 177
R1I3537 N1I353TP1 NVSS 198
R1I3538 N1I353TP5 NVSS 0.21
R1I3539 N1I353TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cioit25s2 DIN E PAD Q
C1I32310 PAD N1I323TP0 235FF
C1I32311 N1I323TP2 PAD 235FF
M1I3230 N1I323TP7 N1I323TP0 NVDD NVDD pch W=38U L=0.34U
M1I3231 N1I323TP0 N1I323TP1 NVDD NVDD pch W=6U L=6U
M1I3232 N1I323TP2 N1I323TP3 NVSS NVSS nch W=6U L=6U
M1I3233 N1I323TP4 N1I323TP2 N1I323TP5 NVSS nch W=38U L=0.34U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E VSS VSS nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=13U L=0.24U
M6 TP2 E TP3 VSS nch W=10U L=0.24U
M7 TP3 TP1 VSS VSS nch W=7.2U L=0.24U
M8 VDD TP20 TP2 VDD pch W=13U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 VSS TP20 TP3 VSS nch W=7.2U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=35.5U L=0.34U
M14 TP14 TP3 NVSS VSS nch W=10.8U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=35.5U L=0.34U
M18 TP15 TP3 NVSS VSS nch W=10.8U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=35.5U L=0.34U
M22 TP16 TP3 NVSS VSS nch W=10.8U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=35.5U L=0.34U
M26 TP17 TP3 NVSS VSS nch W=10.8U L=0.34U
M27 PAD NVSS NVSS VSS nch W=24U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 VSS TP4 Q VSS nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 VSS TP13 TP4 VSS nch W=4.1U L=0.24U
M33 TP20 DIN VDD VDD pch W=3U L=0.24U
M34 TP20 DIN VSS VSS nch W=7U L=0.24U
R1I3234 N1I323TP7 EVSS 123
R1I3235 NVDD N1I323TP3 198
R1I3236 EVDD N1I323TP4 177
R1I3237 N1I323TP1 NVSS 198
R1I3238 N1I323TP5 NVSS 0.21
R1I3239 N1I323TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cioit25s3 DIN E PAD Q
C1I32810 PAD N1I328TP0 235FF
C1I32811 N1I328TP2 PAD 235FF
M1I3280 N1I328TP7 N1I328TP0 NVDD NVDD pch W=38U L=0.34U
M1I3281 N1I328TP0 N1I328TP1 NVDD NVDD pch W=6U L=6U
M1I3282 N1I328TP2 N1I328TP3 NVSS NVSS nch W=6U L=6U
M1I3283 N1I328TP4 N1I328TP2 N1I328TP5 NVSS nch W=38U L=0.34U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E VSS VSS nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=14U L=0.24U
M6 TP2 E TP3 VSS nch W=10U L=0.24U
M7 TP3 TP1 VSS VSS nch W=7.6U L=0.24U
M8 VDD TP20 TP2 VDD pch W=14U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 VSS TP20 TP3 VSS nch W=7.6U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=84U L=0.34U
M14 TP14 TP3 NVSS VSS nch W=24.5U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=84U L=0.34U
M18 TP15 TP3 NVSS VSS nch W=24.5U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=84U L=0.34U
M22 TP16 TP3 NVSS VSS nch W=24.5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=84U L=0.34U
M26 TP17 TP3 NVSS VSS nch W=24.5U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 VSS TP4 Q VSS nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 VSS TP13 TP4 VSS nch W=4.1U L=0.24U
M33 TP20 DIN VDD VDD pch W=3U L=0.24U
M34 TP20 DIN VSS VSS nch W=7U L=0.24U
R1I3284 N1I328TP7 EVSS 123
R1I3285 NVDD N1I328TP3 198
R1I3286 EVDD N1I328TP4 177
R1I3287 N1I328TP1 NVSS 198
R1I3288 N1I328TP5 NVSS 0.21
R1I3289 N1I328TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT cioit25s4 DIN E PAD Q
C1I32410 PAD N1I324TP0 235FF
C1I32411 N1I324TP2 PAD 235FF
M1I3240 N1I324TP7 N1I324TP0 NVDD NVDD pch W=38U L=0.34U
M1I3241 N1I324TP0 N1I324TP1 NVDD NVDD pch W=6U L=6U
M1I3242 N1I324TP2 N1I324TP3 NVSS NVSS nch W=6U L=6U
M1I3243 N1I324TP4 N1I324TP2 N1I324TP5 NVSS nch W=38U L=0.34U
M3 TP20 E VDD VDD pch W=6U L=0.24U
M4 TP20 E VSS VSS nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=18U L=0.24U
M6 TP2 E TP3 VSS nch W=10U L=0.24U
M7 TP3 TP20 VSS VSS nch W=10U L=0.24U
M8 VDD TP1 TP2 VDD pch W=18U L=0.24U
M9 TP2 TP20 TP3 VDD pch W=10U L=0.24U
M10 VSS TP1 TP3 VSS nch W=10U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=152U L=0.34U
M14 TP14 TP3 NVSS VSS nch W=40.8U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=152U L=0.34U
M18 TP15 TP3 NVSS VSS nch W=40.8U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=152U L=0.34U
M22 TP16 TP3 NVSS VSS nch W=40.5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=152U L=0.34U
M26 TP17 TP3 NVSS VSS nch W=40.8U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 VSS TP4 Q VSS nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 VSS TP13 TP4 VSS nch W=4.1U L=0.24U
M33 TP1 DIN VDD VDD pch W=3U L=0.24U
M34 TP1 DIN VSS VSS nch W=7U L=0.24U
R1I3244 N1I324TP7 EVSS 123
R1I3245 NVDD N1I324TP3 198
R1I3246 EVDD N1I324TP4 177
R1I3247 N1I324TP1 NVSS 198
R1I3248 N1I324TP5 NVSS 0.21
R1I3249 N1I324TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ciont25s1 DIN E PAD Q
C1I35310 PAD N1I353TP0 235FF
C1I35311 N1I353TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6U L=0.24U
M1I3530 N1I353TP7 N1I353TP0 NVDD NVDD pch W=38U L=0.34U
M1I3531 N1I353TP0 N1I353TP1 NVDD NVDD pch W=6U L=6U
M1I3532 N1I353TP2 N1I353TP3 NVSS NVSS nch W=6U L=6U
M1I3533 N1I353TP4 N1I353TP2 N1I353TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN VSS VSS nch W=2U L=0.24U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E VSS VSS nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=13U L=0.24U
M6 TP2 E TP3 VSS nch W=10U L=0.24U
M7 TP3 TP1 VSS VSS nch W=7U L=0.24U
M8 VDD TP20 TP2 VDD pch W=13U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 VSS TP20 TP3 VSS nch W=7U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=15.5U L=0.34U
M14 TP14 TP3 NVSS VSS nch W=5U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=15.5U L=0.34U
M18 TP15 TP3 NVSS VSS nch W=5U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=15.5U L=0.34U
M22 TP16 TP3 NVSS VSS nch W=5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=15.5U L=0.34U
M26 TP17 TP3 NVSS VSS nch W=5U L=0.34U
M27 PAD NVSS NVSS VSS nch W=34U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 VSS TP4 Q VSS nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 VSS TP13 TP4 VSS nch W=4.1U L=0.24U
M33 TP20 TP0 VDD VDD pch W=5.4U L=0.24U
M34 TP20 TP0 VSS VSS nch W=7U L=0.24U
R1I3534 N1I353TP7 EVSS 123
R1I3535 NVDD N1I353TP3 198
R1I3536 EVDD N1I353TP4 177
R1I3537 N1I353TP1 NVSS 198
R1I3538 N1I353TP5 NVSS 0.21
R1I3539 N1I353TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ciont25s2 DIN E PAD Q
C1I32310 PAD N1I323TP0 235FF
C1I32311 N1I323TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6U L=0.24U
M1I3230 N1I323TP7 N1I323TP0 NVDD NVDD pch W=38U L=0.34U
M1I3231 N1I323TP0 N1I323TP1 NVDD NVDD pch W=6U L=6U
M1I3232 N1I323TP2 N1I323TP3 NVSS NVSS nch W=6U L=6U
M1I3233 N1I323TP4 N1I323TP2 N1I323TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN VSS VSS nch W=2U L=0.24U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E VSS VSS nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=13U L=0.24U
M6 TP2 E TP3 VSS nch W=10U L=0.24U
M7 TP3 TP1 VSS VSS nch W=7.2U L=0.24U
M8 VDD TP20 TP2 VDD pch W=13U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 VSS TP20 TP3 VSS nch W=7.2U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=35.5U L=0.34U
M14 TP14 TP3 NVSS VSS nch W=10.8U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=35.5U L=0.34U
M18 TP15 TP3 NVSS VSS nch W=10.8U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=35.5U L=0.34U
M22 TP16 TP3 NVSS VSS nch W=10.8U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=35.5U L=0.34U
M26 TP17 TP3 NVSS VSS nch W=10.8U L=0.34U
M27 PAD NVSS NVSS VSS nch W=24U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 VSS TP4 Q VSS nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 VSS TP13 TP4 VSS nch W=4.1U L=0.24U
M33 TP20 TP0 VDD VDD pch W=3U L=0.24U
M34 TP20 TP0 VSS VSS nch W=7U L=0.24U
R1I3234 N1I323TP7 EVSS 123
R1I3235 NVDD N1I323TP3 198
R1I3236 EVDD N1I323TP4 177
R1I3237 N1I323TP1 NVSS 198
R1I3238 N1I323TP5 NVSS 0.21
R1I3239 N1I323TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ciont25s3 DIN E PAD Q
C1I32810 PAD N1I328TP0 235FF
C1I32811 N1I328TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6U L=0.24U
M1I3280 N1I328TP7 N1I328TP0 NVDD NVDD pch W=38U L=0.34U
M1I3281 N1I328TP0 N1I328TP1 NVDD NVDD pch W=6U L=6U
M1I3282 N1I328TP2 N1I328TP3 NVSS NVSS nch W=6U L=6U
M1I3283 N1I328TP4 N1I328TP2 N1I328TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN VSS VSS nch W=2U L=0.24U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E VSS VSS nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=14U L=0.24U
M6 TP2 E TP3 VSS nch W=10U L=0.24U
M7 TP3 TP1 VSS VSS nch W=7.6U L=0.24U
M8 VDD TP20 TP2 VDD pch W=14U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 VSS TP20 TP3 VSS nch W=7.6U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=84U L=0.34U
M14 TP14 TP3 NVSS VSS nch W=24.5U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=84U L=0.34U
M18 TP15 TP3 NVSS VSS nch W=24.5U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=84U L=0.34U
M22 TP16 TP3 NVSS VSS nch W=24.5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=84U L=0.34U
M26 TP17 TP3 NVSS VSS nch W=24.5U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 VSS TP4 Q VSS nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 VSS TP13 TP4 VSS nch W=4.1U L=0.24U
M33 TP20 TP0 VDD VDD pch W=3U L=0.24U
M34 TP20 TP0 VSS VSS nch W=7U L=0.24U
R1I3284 N1I328TP7 EVSS 123
R1I3285 NVDD N1I328TP3 198
R1I3286 EVDD N1I328TP4 177
R1I3287 N1I328TP1 NVSS 198
R1I3288 N1I328TP5 NVSS 0.21
R1I3289 N1I328TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ciont25s4 DIN E PAD Q
C1I32410 PAD N1I324TP0 235FF
C1I32411 N1I324TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6U L=0.24U
M1I3240 N1I324TP7 N1I324TP0 NVDD NVDD pch W=38U L=0.34U
M1I3241 N1I324TP0 N1I324TP1 NVDD NVDD pch W=6U L=6U
M1I3242 N1I324TP2 N1I324TP3 NVSS NVSS nch W=6U L=6U
M1I3243 N1I324TP4 N1I324TP2 N1I324TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN VSS VSS nch W=2U L=0.24U
M3 TP20 E VDD VDD pch W=6U L=0.24U
M4 TP20 E VSS VSS nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=18U L=0.24U
M6 TP2 E TP3 VSS nch W=10U L=0.24U
M7 TP3 TP20 VSS VSS nch W=10U L=0.24U
M8 VDD TP1 TP2 VDD pch W=18U L=0.24U
M9 TP2 TP20 TP3 VDD pch W=10U L=0.24U
M10 VSS TP1 TP3 VSS nch W=10U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=152U L=0.34U
M14 TP14 TP3 NVSS VSS nch W=40.8U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=152U L=0.34U
M18 TP15 TP3 NVSS VSS nch W=40.8U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=152U L=0.34U
M22 TP16 TP3 NVSS VSS nch W=40.5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=152U L=0.34U
M26 TP17 TP3 NVSS VSS nch W=40.8U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 VSS TP4 Q VSS nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 VSS TP13 TP4 VSS nch W=4.1U L=0.24U
M33 TP1 TP0 VDD VDD pch W=3U L=0.24U
M34 TP1 TP0 VSS VSS nch W=7U L=0.24U
R1I3244 N1I324TP7 EVSS 123
R1I3245 NVDD N1I324TP3 198
R1I3246 EVDD N1I324TP4 177
R1I3247 N1I324TP1 NVSS 198
R1I3248 N1I324TP5 NVSS 0.21
R1I3249 N1I324TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT coi25s1 DIN PAD
C1I46610 PAD N1I466TP0 235FF
C1I46611 N1I466TP2 PAD 235FF
M1I4660 N1I466TP7 N1I466TP0 NVDD NVDD pch W=38U L=0.34U
M1I4661 N1I466TP0 N1I466TP1 NVDD NVDD pch W=6U L=6U
M1I4662 N1I466TP2 N1I466TP3 NVSS NVSS nch W=6U L=6U
M1I4663 N1I466TP4 N1I466TP2 N1I466TP5 NVSS nch W=38U L=0.34U
M3 TP1 DIN VDD VDD pch W=7.3U L=0.24U
M4 TP1 DIN VSS VSS nch W=5.2U L=0.24U
M5 TP2 TP1 VDD VDD pch W=23.3U L=0.24U
M6 TP2 TP1 VSS VSS nch W=9.2U L=0.24U
M7 TP3 TP2 NVDD VDD pch W=19U L=0.34U
M8 TP7 TP2 NVSS VSS nch W=6.5U L=0.34U
M9 TP4 TP2 NVDD VDD pch W=19U L=0.34U
M10 TP8 TP2 NVSS VSS nch W=6.5U L=0.34U
M11 TP5 TP2 NVDD VDD pch W=19U L=0.34U
M12 TP9 TP2 NVSS VSS nch W=6.5U L=0.34U
M13 TP6 TP2 NVDD VDD pch W=19U L=0.34U
M14 TP10 TP2 NVSS VSS nch W=6.5U L=0.34U
M15 PAD NVSS NVSS VSS nch W=20U L=0.34U
R1I4664 N1I466TP7 EVSS 123
R1I4665 NVDD N1I466TP3 198
R1I4666 EVDD N1I466TP4 177
R1I4667 N1I466TP1 NVSS 198
R1I4668 N1I466TP5 NVSS 0.21
R1I4669 N1I466TP5 NVSS 0.21
R15 TP3 PAD 17
R16 TP4 PAD 17
R17 TP5 PAD 17
R18 TP6 PAD 17
R19 PAD TP7 17
R20 PAD TP8 17
R21 PAD TP9 17
R22 PAD TP10 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT coi25s4 DIN PAD
C1I44310 PAD N1I443TP0 235FF
C1I44311 N1I443TP2 PAD 235FF
M1I4430 N1I443TP7 N1I443TP0 NVDD NVDD pch W=38U L=0.34U
M1I4431 N1I443TP0 N1I443TP1 NVDD NVDD pch W=6U L=6U
M1I4432 N1I443TP2 N1I443TP3 NVSS NVSS nch W=6U L=6U
M1I4433 N1I443TP4 N1I443TP2 N1I443TP5 NVSS nch W=38U L=0.34U
M3 TP1 DIN VDD VDD pch W=9.3U L=0.24U
M4 TP1 DIN VSS VSS nch W=6.4U L=0.24U
M5 TP2 TP1 VDD VDD pch W=42.1U L=0.24U
M6 TP2 TP1 VSS VSS nch W=17.2U L=0.24U
M7 TP3 TP2 NVDD VDD pch W=124U L=0.34U
M8 TP34 TP2 NVSS VSS nch W=40.5U L=0.34U
M9 TP31 TP2 NVDD VDD pch W=124U L=0.34U
M10 TP35 TP2 NVSS VSS nch W=40.5U L=0.34U
M11 TP32 TP2 NVDD VDD pch W=124U L=0.34U
M12 TP36 TP2 NVSS VSS nch W=40.5U L=0.34U
M13 TP33 TP2 NVDD VDD pch W=124U L=0.34U
M14 TP37 TP2 NVSS VSS nch W=40.5U L=0.34U
R1I4434 N1I443TP7 EVSS 123
R1I4435 NVDD N1I443TP3 198
R1I4436 EVDD N1I443TP4 177
R1I4437 N1I443TP1 NVSS 198
R1I4438 N1I443TP5 NVSS 0.21
R1I4439 N1I443TP5 NVSS 0.21
R15 TP3 PAD 17
R16 TP31 PAD 17
R17 TP32 PAD 17
R18 TP33 PAD 17
R19 PAD TP34 17
R20 PAD TP35 17
R21 PAD TP36 17
R22 PAD TP37 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT con25s1 DIN PAD
C1I46710 PAD N1I467TP0 235FF
C1I46711 N1I467TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6.2U L=0.24U
M1I4670 N1I467TP7 N1I467TP0 NVDD NVDD pch W=38U L=0.34U
M1I4671 N1I467TP0 N1I467TP1 NVDD NVDD pch W=6U L=6U
M1I4672 N1I467TP2 N1I467TP3 NVSS NVSS nch W=6U L=6U
M1I4673 N1I467TP4 N1I467TP2 N1I467TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN VSS VSS nch W=3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=7.3U L=0.24U
M4 TP1 TP0 VSS VSS nch W=5.2U L=0.24U
M5 TP2 TP1 VDD VDD pch W=23.3U L=0.24U
M6 TP2 TP1 VSS VSS nch W=9.2U L=0.24U
M7 TP3 TP2 NVDD VDD pch W=19U L=0.34U
M8 TP7 TP2 NVSS VSS nch W=6.5U L=0.34U
M9 TP4 TP2 NVDD VDD pch W=19U L=0.34U
M10 TP8 TP2 NVSS VSS nch W=6.5U L=0.34U
M11 TP5 TP2 NVDD VDD pch W=19U L=0.34U
M12 TP9 TP2 NVSS VSS nch W=6.5U L=0.34U
M13 TP6 TP2 NVDD VDD pch W=19U L=0.34U
M14 TP10 TP2 NVSS VSS nch W=6.5U L=0.34U
M15 PAD NVSS NVSS VSS nch W=20U L=0.34U
R1I4674 N1I467TP7 EVSS 123
R1I4675 NVDD N1I467TP3 198
R1I4676 EVDD N1I467TP4 177
R1I4677 N1I467TP1 NVSS 198
R1I4678 N1I467TP5 NVSS 0.21
R1I4679 N1I467TP5 NVSS 0.21
R15 TP3 PAD 17
R16 TP4 PAD 17
R17 TP5 PAD 17
R18 TP6 PAD 17
R19 PAD TP7 17
R20 PAD TP8 17
R21 PAD TP9 17
R22 PAD TP10 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT con25s4 DIN PAD
C1I44410 PAD N1I444TP0 235FF
C1I44411 N1I444TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6.2U L=0.24U
M1I4440 N1I444TP7 N1I444TP0 NVDD NVDD pch W=38U L=0.34U
M1I4441 N1I444TP0 N1I444TP1 NVDD NVDD pch W=6U L=6U
M1I4442 N1I444TP2 N1I444TP3 NVSS NVSS nch W=6U L=6U
M1I4443 N1I444TP4 N1I444TP2 N1I444TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN VSS VSS nch W=3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=9.3U L=0.24U
M4 TP1 TP0 VSS VSS nch W=6.4U L=0.24U
M5 TP2 TP1 VDD VDD pch W=42.1U L=0.24U
M6 TP2 TP1 VSS VSS nch W=17.2U L=0.24U
M7 TP3 TP2 NVDD VDD pch W=124U L=0.34U
M8 TP34 TP2 NVSS VSS nch W=40.5U L=0.34U
M9 TP31 TP2 NVDD VDD pch W=124U L=0.34U
M10 TP35 TP2 NVSS VSS nch W=40.5U L=0.34U
M11 TP32 TP2 NVDD VDD pch W=124U L=0.34U
M12 TP36 TP2 NVSS VSS nch W=40.5U L=0.34U
M13 TP33 TP2 NVDD VDD pch W=124U L=0.34U
M14 TP37 TP2 NVSS VSS nch W=40.5U L=0.34U
R1I4444 N1I444TP7 EVSS 123
R1I4445 NVDD N1I444TP3 198
R1I4446 EVDD N1I444TP4 177
R1I4447 N1I444TP1 NVSS 198
R1I4448 N1I444TP5 NVSS 0.21
R1I4449 N1I444TP5 NVSS 0.21
R15 TP3 PAD 17
R16 TP31 PAD 17
R17 TP32 PAD 17
R18 TP33 PAD 17
R19 PAD TP34 17
R20 PAD TP35 17
R21 PAD TP36 17
R22 PAD TP37 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT corner INOUT2 INOUT1 AVCC AVSS VCC VSS NVCC NVSS
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ncdavdd NVDD VDD AVDD EVDD PAD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 EVDD N1N43 NVSS NVSS nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N43 NVSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 NVDD PAD 0.0003
R3 AVDD VDD 0.0016
R4 VDD NVDD 0.0016
R5 EVDD PAD 0.0016
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ncdavss NVSS VSS AVSS EVSS PAD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 EVSS N1N85 NVDD NVDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 NVDD N1N85 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 EVSS PAD 0.0024
R3 NVSS PAD 0.000966
R4 AVSS VSS 0.002
R5 VSS EVSS 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ncdvdd NVDD PAD VDD EVDD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 EVDD N1N43 NVSS NVSS nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N43 NVSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 NVDD PAD 0.003
R3 NVDD VDD 0.0016
R4 PAD EVDD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ncdvss NVSS PAD VSS EVSS
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 VSS N1N85 NVDD NVDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 NVDD N1N85 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 EVSS PAD 0.002
R3 NVSS PAD 0.002
R4 VSS EVSS 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ndavdd NVDD PAD AVDD EVDD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 EVDD N1N44 NVSS NVSS nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N44 NVSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 NVDD PAD 0.002
R3 AVDD NVDD 0.002
R4 EVDD PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ndavss NVSS PAD EVSS AVSS
C1I6210 PAD N1I62TP0 235FF
C1I6211 N1I62TP2 PAD 235FF
M1 EVSS N1N56 NVDD NVDD pch W=300U L=0.34U
M1I620 N1I62TP7 N1I62TP0 NVDD NVDD pch W=38U L=0.34U
M1I621 N1I62TP0 N1I62TP1 NVDD NVDD pch W=6U L=6U
M1I622 N1I62TP2 N1I62TP3 NVSS NVSS nch W=6U L=6U
M1I623 N1I62TP4 N1I62TP2 N1I62TP5 NVSS nch W=38U L=0.34U
R1 NVDD N1N56 400
R1I624 N1I62TP7 EVSS 123
R1I625 NVDD N1I62TP3 198
R1I626 EVDD N1I62TP4 177
R1I627 N1I62TP1 NVSS 198
R1I628 N1I62TP5 NVSS 0.21
R1I629 N1I62TP5 NVSS 0.21
R2 EVSS PAD 0.001
R3 NVSS PAD 0.00035
R4 AVSS EVSS 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ndvdd EVDD NVDD PAD N1
C1I6210 PAD N1I62TP0 235FF
C1I6211 N1I62TP2 PAD 235FF
M1 EVDD N1N44 NVSS NVSS nch W=300U L=0.34U
M1I620 N1I62TP7 N1I62TP0 NVDD NVDD pch W=38U L=0.34U
M1I621 N1I62TP0 N1I62TP1 NVDD NVDD pch W=6U L=6U
M1I622 N1I62TP2 N1I62TP3 NVSS NVSS nch W=6U L=6U
M1I623 N1I62TP4 N1I62TP2 N1I62TP5 NVSS nch W=38U L=0.34U
R1 N1N44 NVSS 400
R1I624 N1I62TP7 EVSS 123
R1I625 NVDD N1I62TP3 198
R1I626 EVDD N1I62TP4 177
R1I627 N1I62TP1 NVSS 198
R1I628 N1I62TP5 NVSS 0.21
R1I629 N1I62TP5 NVSS 0.21
R2 NVDD PAD 0.0023
R3 PAD EVDD 0.0018
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT ndvss NVSS PAD EVSS N1
C1I6210 PAD N1I62TP0 235FF
C1I6211 N1I62TP2 PAD 235FF
M1 EVSS N1N56 NVDD NVDD pch W=300U L=0.34U
M1I620 N1I62TP7 N1I62TP0 NVDD NVDD pch W=38U L=0.34U
M1I621 N1I62TP0 N1I62TP1 NVDD NVDD pch W=6U L=6U
M1I622 N1I62TP2 N1I62TP3 NVSS NVSS nch W=6U L=6U
M1I623 N1I62TP4 N1I62TP2 N1I62TP5 NVSS nch W=38U L=0.34U
R1 NVDD N1N56 400
R1I624 N1I62TP7 EVSS 123
R1I625 NVDD N1I62TP3 198
R1I626 EVDD N1I62TP4 177
R1I627 N1I62TP1 NVSS 198
R1I628 N1I62TP5 NVSS 0.21
R1I629 N1I62TP5 NVSS 0.21
R2 NVSS PAD 0.0027
R3 EVSS PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and2s1 Q DIN1 DIN2
M1 N1N251 DIN1 VDD VDD pch W=0.7U L=0.24U
M2 N1N251 DIN2 VDD VDD pch W=0.7U L=0.24U
M3 N1N251 DIN1 N1N257 0 nch W=0.7U L=0.24U
M4 N1N257 DIN2 GVSS 0 nch W=0.7U L=0.24U
M5 Q N1N251 VDD VDD pch W=1.76U L=0.24U
M6 Q N1N251 GVSS 0 nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and2s2 Q DIN1 DIN2
M3 N1N257 DIN1 N1N259 0 nch W=2.14U L=0.24U
M1 N1N257 DIN1 VDD VDD pch W=2.4U L=0.24U
M2 N1N257 DIN2 VDD VDD pch W=2.4U L=0.24U
M5 Q N1N257 VDD VDD pch W=5.3U L=0.24U
M4 N1N259 DIN2 GVSS 0 nch W=2.14U L=0.24U
M6 Q N1N257 GVSS 0 nch W=3.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and2s3 Q DIN1 DIN2
M3 N1N257 DIN1 N1N259 0 nch W=4.4U L=0.24U
M1 N1N257 DIN1 VDD VDD pch W=4.5U L=0.24U
M2 N1N257 DIN2 VDD VDD pch W=4.5U L=0.24U
M4 N1N259 DIN2 GVSS 0 nch W=4.4U L=0.24U
M5 Q N1N257 VDD VDD pch W=9.5U L=0.24U
M6 Q N1N257 GVSS 0 nch W=6.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and3s1 Q DIN1 DIN2 DIN3
M4 N1N258 DIN1 N1N262 0 nch W=1.08U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=0.82U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=0.82U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=0.82U L=0.24U
M5 N1N262 DIN2 N1N264 0 nch W=1.08U L=0.24U
M6 N1N264 DIN3 GVSS 0 nch W=1.08U L=0.24U
M8 Q N1N258 GVSS 0 nch W=1.34U L=0.24U
M7 Q N1N258 VDD VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and3s2 Q DIN1 DIN2 DIN3
M4 N1N258 DIN1 N1N262 0 nch W=3.14U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=2.54U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=2.54U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=2.54U L=0.24U
M5 N1N262 DIN2 N1N264 0 nch W=3.14U L=0.24U
M6 N1N264 DIN3 GVSS 0 nch W=3.14U L=0.24U
M8 Q N1N258 GVSS 0 nch W=4.1U L=0.24U
M7 Q N1N258 VDD VDD pch W=4.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and3s3 Q DIN1 DIN2 DIN3
M4 N1N258 DIN1 N1N262 0 nch W=3.8U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=4.7U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=4.7U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=4.7U L=0.24U
M5 N1N262 DIN2 N1N264 0 nch W=4.76U L=0.24U
M6 N1N264 DIN3 GVSS 0 nch W=7.4U L=0.24U
M8 Q N1N258 GVSS 0 nch W=7.4U L=0.24U
M7 Q N1N258 VDD VDD pch W=9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and4s1 Q DIN1 DIN2 DIN3 DIN4
M5 N1N258 DIN1 N1N265 0 nch W=1U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=1U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=1U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=1U L=0.24U
M4 N1N258 DIN4 VDD VDD pch W=1U L=0.24U
M6 N1N265 DIN2 N1N267 0 nch W=1.24U L=0.24U
M7 N1N267 DIN3 N1N269 0 nch W=1.44U L=0.24U
M8 N1N269 DIN4 GVSS 0 nch W=1.64U L=0.24U
M9 Q N1N258 VDD VDD pch W=1.96U L=0.24U
M10 Q N1N258 GVSS 0 nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and4s2 Q DIN1 DIN2 DIN3 DIN4
M5 N1N258 DIN1 N1N265 0 nch W=2.32U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=3U L=0.24U
M2 N1N258 DIN2 VDD VDD pch W=3U L=0.24U
M3 N1N258 DIN3 VDD VDD pch W=3U L=0.24U
M4 N1N258 DIN4 VDD VDD pch W=3U L=0.24U
M6 N1N265 DIN2 N1N267 0 nch W=2.54U L=0.24U
M7 N1N267 DIN3 N1N269 0 nch W=3.96U L=0.24U
M8 N1N269 DIN4 GVSS 0 nch W=4.16U L=0.24U
M9 Q N1N258 VDD VDD pch W=5.7U L=0.24U
M10 Q N1N258 GVSS 0 nch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_and4s3 DIN1 DIN2 DIN3 DIN4 Q
M3 N1N259 DIN1 N1N262 0 nch W=3.16U L=0.24U
M1 N1N259 DIN1 VDD VDD pch W=3.5U L=0.24U
M2 VDD DIN2 N1N259 VDD pch W=3.5U L=0.24U
M4 N1N262 DIN2 GVSS 0 nch W=4.1U L=0.24U
M9 N1N279 N1N259 VDD VDD pch W=7.2U L=0.24U
M10 N1N279 N1N270 Q VDD pch W=7U L=0.24U
M5 N1N270 DIN3 VDD VDD pch W=3.5U L=0.24U
M6 VDD DIN4 N1N270 VDD pch W=3.5U L=0.24U
M7 N1N270 DIN3 N1N273 0 nch W=3.16U L=0.24U
M8 N1N273 DIN4 GVSS 0 nch W=4.1U L=0.24U
M11 Q N1N259 GVSS 0 nch W=2.5U L=0.24U
M12 GVSS N1N270 Q 0 nch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoai1112s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N286 DIN1 Q 0 nch W=0.8U L=0.24U
M1 N1N282 DIN4 VDD VDD pch W=1.5U L=0.24U
M2 N1N282 DIN5 VDD VDD pch W=1.5U L=0.24U
M3 Q DIN3 N1N282 VDD pch W=1.4U L=0.24U
M4 VDD DIN2 Q VDD pch W=0.7U L=0.24U
M5 VDD DIN1 Q VDD pch W=0.7U L=0.24U
M7 N1N299 DIN2 N1N286 0 nch W=0.8U L=0.24U
M8 N1N299 DIN3 GVSS 0 nch W=0.8U L=0.24U
M9 N1N299 DIN4 N1N302 0 nch W=1.6U L=0.24U
M10 N1N302 DIN5 GVSS 0 nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoai1112s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N286 DIN1 Q 0 nch W=1.1U L=0.24U
M1 N1N282 DIN4 VDD VDD pch W=2U L=0.24U
M2 N1N282 DIN5 VDD VDD pch W=2U L=0.24U
M3 Q DIN3 N1N282 VDD pch W=1.9U L=0.24U
M4 VDD DIN2 Q VDD pch W=1U L=0.24U
M5 VDD DIN1 Q VDD pch W=1U L=0.24U
M7 N1N299 DIN2 N1N286 0 nch W=1.1U L=0.24U
M8 N1N299 DIN3 GVSS 0 nch W=1.1U L=0.24U
M9 N1N299 DIN4 N1N302 0 nch W=2.2U L=0.24U
M10 N1N302 DIN5 GVSS 0 nch W=2.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoai1112s3 DIN1 DIN2 DIN3 DIN4 DIN5 Q
M6 N1N286 DIN1 Q 0 nch W=1.6U L=0.24U
M1 N1N282 DIN4 VDD VDD pch W=3.3U L=0.24U
M2 N1N282 DIN5 VDD VDD pch W=3.4U L=0.24U
M3 Q DIN3 N1N282 VDD pch W=3.3U L=0.24U
M4 VDD DIN2 Q VDD pch W=1.7U L=0.24U
M5 VDD DIN1 Q VDD pch W=1.7U L=0.24U
M7 N1N299 DIN2 N1N286 0 nch W=1.7U L=0.24U
M8 N1N299 DIN3 GVSS 0 nch W=1.7U L=0.24U
M9 N1N299 DIN4 N1N302 0 nch W=3.4U L=0.24U
M10 N1N302 DIN5 GVSS 0 nch W=3.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoai122s1 DIN1 DIN2 DIN3 DIN4 DIN5 Q
M6 Q DIN1 N1N298 0 nch W=0.9U L=0.24U
M2 N1N290 DIN2 VDD VDD pch W=1.5U L=0.24U
M3 Q DIN4 N1N290 VDD pch W=1.5U L=0.24U
M4 VDD DIN3 N1N290 VDD pch W=1.5U L=0.24U
M5 N1N290 DIN5 Q VDD pch W=1.5U L=0.24U
M7 N1N298 DIN2 N1N300 0 nch W=0.9U L=0.24U
M10 GVSS DIN5 N1N302 0 nch W=0.9U L=0.24U
M9 N1N302 DIN4 N1N298 0 nch W=0.9U L=0.24U
M8 GVSS DIN3 N1N300 0 nch W=0.9U L=0.24U
M1 Q DIN1 VDD VDD pch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoai122s2 DIN1 DIN2 DIN3 DIN4 DIN5 Q
M6 Q DIN1 N1N298 0 nch W=1.1U L=0.24U
M2 N1N290 DIN2 VDD VDD pch W=1.8U L=0.24U
M3 Q DIN4 N1N290 VDD pch W=1.8U L=0.24U
M4 VDD DIN3 N1N290 VDD pch W=1.8U L=0.24U
M5 N1N290 DIN5 Q VDD pch W=1.8U L=0.24U
M7 N1N298 DIN2 N1N300 0 nch W=1.1U L=0.24U
M10 GVSS DIN5 N1N302 0 nch W=1.1U L=0.24U
M9 N1N302 DIN4 N1N298 0 nch W=1.1U L=0.24U
M8 GVSS DIN3 N1N300 0 nch W=1.1U L=0.24U
M1 Q DIN1 VDD VDD pch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoai122s3 DIN1 DIN2 DIN3 DIN4 DIN5 Q
M6 N1N292 DIN1 N1N298 0 nch W=0.9U L=0.24U
M2 N1N290 DIN2 VDD VDD pch W=1.5U L=0.24U
M3 N1N292 DIN4 N1N290 VDD pch W=1.5U L=0.24U
M4 VDD DIN3 N1N290 VDD pch W=1.5U L=0.24U
M5 N1N290 DIN5 N1N292 VDD pch W=1.5U L=0.24U
M7 N1N298 DIN2 N1N300 0 nch W=1U L=0.24U
M10 GVSS DIN5 N1N302 0 nch W=1U L=0.24U
M9 N1N302 DIN4 N1N298 0 nch W=1U L=0.24U
M8 GVSS DIN3 N1N300 0 nch W=1U L=0.24U
M1 N1N292 DIN1 VDD VDD pch W=0.7U L=0.24U
M12 N1N339 N1N292 GVSS 0 nch W=1.4U L=0.24U
M11 N1N339 N1N292 VDD VDD pch W=2.7U L=0.24U
M13 Q N1N339 VDD VDD pch W=4.5U L=0.24U
M14 Q N1N339 GVSS 0 nch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi123s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N461 DIN3 N1N445 VDD pch W=4.1U L=0.24U
M1 N1N445 DIN5 VDD VDD pch W=4.1U L=0.24U
M2 VDD DIN4 N1N445 VDD pch W=4.1U L=0.24U
M3 VDD DIN6 N1N445 VDD pch W=4.1U L=0.24U
M5 N1N445 DIN2 N1N461 VDD pch W=4.1U L=0.24U
M6 Q DIN1 N1N461 VDD pch W=4.1U L=0.24U
M7 N1N469 DIN2 Q 0 nch W=1.2U L=0.24U
M10 N1N469 DIN3 GVSS 0 nch W=1.2U L=0.24U
M8 N1N473 DIN4 Q 0 nch W=1.8U L=0.24U
M12 GVSS DIN6 N1N475 0 nch W=1.8U L=0.24U
M11 N1N475 DIN5 N1N473 0 nch W=1.8U L=0.24U
M9 Q DIN1 GVSS 0 nch W=0.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi123s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N461 DIN3 N1N445 VDD pch W=5.8U L=0.24U
M1 N1N445 DIN5 VDD VDD pch W=5.8U L=0.24U
M2 VDD DIN4 N1N445 VDD pch W=5.8U L=0.24U
M3 VDD DIN6 N1N445 VDD pch W=5.8U L=0.24U
M5 N1N445 DIN2 N1N461 VDD pch W=5.8U L=0.24U
M6 Q DIN1 N1N461 VDD pch W=5.8U L=0.24U
M7 N1N469 DIN2 Q 0 nch W=1.7U L=0.24U
M10 N1N469 DIN3 GVSS 0 nch W=1.7U L=0.24U
M8 N1N473 DIN4 Q 0 nch W=2.5U L=0.24U
M12 GVSS DIN6 N1N475 0 nch W=2.5U L=0.24U
M11 N1N475 DIN5 N1N473 0 nch W=2.5U L=0.24U
M9 Q DIN1 GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi123s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N461 DIN3 N1N445 VDD pch W=7.8U L=0.24U
M1 N1N445 DIN5 VDD VDD pch W=7.8U L=0.24U
M2 VDD DIN4 N1N445 VDD pch W=7.8U L=0.24U
M3 VDD DIN6 N1N445 VDD pch W=7.8U L=0.24U
M5 N1N445 DIN2 N1N461 VDD pch W=7.8U L=0.24U
M6 Q DIN1 N1N461 VDD pch W=7.8U L=0.24U
M7 N1N469 DIN2 Q 0 nch W=2.2U L=0.24U
M10 N1N469 DIN3 GVSS 0 nch W=2.2U L=0.24U
M8 N1N473 DIN4 Q 0 nch W=3.3U L=0.24U
M12 GVSS DIN6 N1N475 0 nch W=3.3U L=0.24U
M11 N1N475 DIN5 N1N473 0 nch W=3.3U L=0.24U
M9 Q DIN1 GVSS 0 nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi13s1 Q DIN1 DIN2 DIN3 DIN4
M6 N1N452 DIN2 Q 0 nch W=1.24U L=0.24U
M2 VDD DIN3 N1N490 VDD pch W=2.8U L=0.24U
M5 Q DIN1 GVSS 0 nch W=0.6U L=0.24U
M4 Q DIN1 N1N490 VDD pch W=2.7U L=0.24U
M1 N1N490 DIN2 VDD VDD pch W=2.8U L=0.24U
M3 VDD DIN4 N1N490 VDD pch W=2.8U L=0.24U
M8 GVSS DIN4 N1N454 0 nch W=1U L=0.24U
M7 N1N454 DIN3 N1N452 0 nch W=1.24U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi13s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 GVSS 0 nch W=0.8U L=0.24U
M4 Q DIN1 N1N486 VDD pch W=4U L=0.24U
M1 N1N486 DIN2 VDD VDD pch W=4.1U L=0.24U
M2 VDD DIN3 N1N486 VDD pch W=4.1U L=0.24U
M3 VDD DIN4 N1N486 VDD pch W=4.1U L=0.24U
M6 N1N452 DIN2 Q 0 nch W=1.84U L=0.24U
M7 N1N454 DIN3 N1N452 0 nch W=1.84U L=0.24U
M8 GVSS DIN4 N1N454 0 nch W=1.84U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi13s3 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 GVSS 0 nch W=1U L=0.24U
M4 Q DIN1 N1N486 VDD pch W=6U L=0.24U
M1 N1N486 DIN2 VDD VDD pch W=6U L=0.24U
M2 VDD DIN3 N1N486 VDD pch W=6U L=0.24U
M3 VDD DIN4 N1N486 VDD pch W=6U L=0.24U
M6 N1N452 DIN2 Q 0 nch W=2.8U L=0.24U
M7 N1N454 DIN3 N1N452 0 nch W=2.8U L=0.24U
M8 GVSS DIN4 N1N454 0 nch W=2.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi211s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N444 0 nch W=1U L=0.24U
M3 N1N439 DIN4 N1N477 VDD pch W=3.7U L=0.24U
M4 Q DIN3 N1N477 VDD pch W=3.7U L=0.24U
M2 VDD DIN2 N1N439 VDD pch W=3.8U L=0.24U
M1 N1N439 DIN1 VDD VDD pch W=3.8U L=0.24U
M7 Q DIN3 GVSS 0 nch W=0.6U L=0.24U
M8 GVSS DIN4 Q 0 nch W=0.6U L=0.24U
M6 N1N444 DIN2 GVSS 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi211s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N444 0 nch W=1.3U L=0.24U
M3 N1N439 DIN4 N1N477 VDD pch W=4.8U L=0.24U
M4 Q DIN3 N1N477 VDD pch W=4.7U L=0.24U
M2 VDD DIN2 N1N439 VDD pch W=4.9U L=0.24U
M1 N1N439 DIN1 VDD VDD pch W=4.9U L=0.24U
M7 Q DIN3 GVSS 0 nch W=0.8U L=0.24U
M8 GVSS DIN4 Q 0 nch W=0.8U L=0.24U
M6 N1N444 DIN2 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi211s3 Q DIN1 DIN2 DIN3 DIN4
M5 N1N467 DIN1 N1N444 0 nch W=1.4U L=0.24U
M3 N1N439 DIN4 N1N480 VDD pch W=4.1U L=0.24U
M4 N1N467 DIN3 N1N480 VDD pch W=3.9U L=0.24U
M2 VDD DIN2 N1N439 VDD pch W=4.3U L=0.24U
M1 N1N439 DIN1 VDD VDD pch W=4.3U L=0.24U
M7 N1N467 DIN3 GVSS 0 nch W=0.7U L=0.24U
M8 GVSS DIN4 N1N467 0 nch W=0.7U L=0.24U
M6 N1N444 DIN2 GVSS 0 nch W=1.4U L=0.24U
M9 N1N489 N1N467 VDD VDD pch W=2.4U L=0.24U
M10 N1N489 N1N467 GVSS 0 nch W=1.6U L=0.24U
M12 Q N1N489 GVSS 0 nch W=2U L=0.24U
M11 Q N1N489 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi21s1 Q DIN1 DIN2 DIN3
M5 Q DIN3 GVSS 0 nch W=0.6U L=0.24U
M2 VDD DIN1 N1N344 VDD pch W=2.76U L=0.24U
M3 Q DIN3 N1N344 VDD pch W=2.76U L=0.24U
M1 N1N344 DIN2 VDD VDD pch W=2.76U L=0.24U
M4 Q DIN2 N1N322 0 nch W=1U L=0.24U
M6 N1N322 DIN1 GVSS 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi21s2 Q DIN1 DIN2 DIN3
M5 Q DIN3 GVSS 0 nch W=0.8U L=0.24U
M2 VDD DIN1 N1N344 VDD pch W=3.54U L=0.24U
M3 Q DIN3 N1N344 VDD pch W=3.54U L=0.24U
M1 N1N344 DIN2 VDD VDD pch W=3.54U L=0.24U
M4 Q DIN2 N1N322 0 nch W=1.3U L=0.24U
M6 N1N322 DIN1 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi21s3 Q DIN1 DIN2 DIN3
M5 Q DIN3 GVSS 0 nch W=1U L=0.24U
M2 VDD DIN1 N1N344 VDD pch W=4.6U L=0.24U
M3 Q DIN3 N1N344 VDD pch W=4.6U L=0.24U
M1 N1N344 DIN2 VDD VDD pch W=4.6U L=0.24U
M4 Q DIN2 N1N322 0 nch W=1.7U L=0.24U
M6 N1N322 DIN1 GVSS 0 nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi221s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N449 0 nch W=1U L=0.24U
M1 N1N439 DIN3 VDD VDD pch W=3.6U L=0.24U
M2 VDD DIN4 N1N439 VDD pch W=3.6U L=0.24U
M4 N1N439 DIN2 N1N443 VDD pch W=3.5U L=0.24U
M3 N1N443 DIN1 N1N439 VDD pch W=3.5U L=0.24U
M5 Q DIN5 N1N443 VDD pch W=3.4U L=0.24U
M8 N1N451 DIN3 Q 0 nch W=1U L=0.24U
M10 GVSS DIN4 N1N451 0 nch W=1U L=0.24U
M9 N1N449 DIN2 GVSS 0 nch W=1U L=0.24U
M7 Q DIN5 GVSS 0 nch W=0.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi221s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N449 0 nch W=1.22U L=0.24U
M1 N1N439 DIN3 VDD VDD pch W=4.3U L=0.24U
M3 N1N443 DIN1 N1N439 VDD pch W=4.2U L=0.24U
M5 Q DIN5 N1N443 VDD pch W=4.1U L=0.24U
M2 VDD DIN4 N1N439 VDD pch W=4.3U L=0.24U
M4 N1N439 DIN2 N1N443 VDD pch W=4.2U L=0.24U
M9 N1N449 DIN2 GVSS 0 nch W=1.22U L=0.24U
M7 Q DIN5 GVSS 0 nch W=0.74U L=0.24U
M8 N1N451 DIN3 Q 0 nch W=1.22U L=0.24U
M10 GVSS DIN4 N1N451 0 nch W=1.22U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi221s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N446 DIN1 N1N449 0 nch W=1.3U L=0.24U
M1 N1N439 DIN3 VDD VDD pch W=3.7U L=0.24U
M3 N1N443 DIN1 N1N439 VDD pch W=3.5U L=0.24U
M5 N1N446 DIN5 N1N443 VDD pch W=3.4U L=0.24U
M2 VDD DIN4 N1N439 VDD pch W=3.7U L=0.24U
M4 N1N439 DIN2 N1N443 VDD pch W=3.5U L=0.24U
M9 N1N449 DIN2 GVSS 0 nch W=1.3U L=0.24U
M7 N1N446 DIN5 GVSS 0 nch W=0.7U L=0.24U
M8 N1N451 DIN3 N1N446 0 nch W=1.3U L=0.24U
M10 GVSS DIN4 N1N451 0 nch W=1.3U L=0.24U
M11 N1N527 N1N446 VDD VDD pch W=2.5U L=0.24U
M12 N1N527 N1N446 GVSS 0 nch W=1.6U L=0.24U
M14 Q N1N527 GVSS 0 nch W=2U L=0.24U
M13 Q N1N527 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi2221s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M1 N1N487 DIN1 VDD VDD pch W=5.8U L=0.24U
M3 N1N489 DIN3 N1N487 VDD pch W=5.6U L=0.24U
M5 N1N452 DIN5 N1N489 VDD pch W=5.4U L=0.24U
M2 VDD DIN2 N1N487 VDD pch W=5.8U L=0.24U
M4 N1N487 DIN4 N1N489 VDD pch W=5.6U L=0.24U
M6 N1N489 DIN6 N1N452 VDD pch W=5.4U L=0.24U
M8 Q DIN1 N1N454 0 nch W=1.2U L=0.24U
M9 Q DIN3 N1N506 0 nch W=1.2U L=0.24U
M13 N1N506 DIN4 GVSS 0 nch W=1.2U L=0.24U
M12 N1N454 DIN2 GVSS 0 nch W=1.2U L=0.24U
M10 N1N508 DIN5 Q 0 nch W=1.2U L=0.24U
M14 GVSS DIN6 N1N508 0 nch W=1.2U L=0.24U
M11 GVSS DIN7 Q 0 nch W=0.6U L=0.24U
M7 Q DIN7 N1N452 VDD pch W=5.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi2221s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M1 N1N487 DIN1 VDD VDD pch W=7.1U L=0.24U
M3 N1N489 DIN3 N1N487 VDD pch W=6.9U L=0.24U
M5 N1N452 DIN5 N1N489 VDD pch W=6.7U L=0.24U
M2 VDD DIN2 N1N487 VDD pch W=7.1U L=0.24U
M4 N1N487 DIN4 N1N489 VDD pch W=6.9U L=0.24U
M6 N1N489 DIN6 N1N452 VDD pch W=6.7U L=0.24U
M8 Q DIN1 N1N454 0 nch W=1.4U L=0.24U
M9 Q DIN3 N1N506 0 nch W=1.4U L=0.24U
M13 N1N506 DIN4 GVSS 0 nch W=1.4U L=0.24U
M12 N1N454 DIN2 GVSS 0 nch W=1.4U L=0.24U
M10 N1N508 DIN5 Q 0 nch W=1.4U L=0.24U
M14 GVSS DIN6 N1N508 0 nch W=1.4U L=0.24U
M11 GVSS DIN7 Q 0 nch W=0.7U L=0.24U
M7 Q DIN7 N1N452 VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi2221s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M1 N1N487 DIN1 VDD VDD pch W=8.6U L=0.24U
M3 N1N489 DIN3 N1N487 VDD pch W=8.4U L=0.24U
M5 N1N452 DIN5 N1N489 VDD pch W=8.2U L=0.24U
M2 VDD DIN2 N1N487 VDD pch W=8.6U L=0.24U
M4 N1N487 DIN4 N1N489 VDD pch W=8.4U L=0.24U
M6 N1N489 DIN6 N1N452 VDD pch W=8.2U L=0.24U
M8 Q DIN1 N1N454 0 nch W=1.8U L=0.24U
M9 Q DIN3 N1N506 0 nch W=1.8U L=0.24U
M13 N1N506 DIN4 GVSS 0 nch W=1.8U L=0.24U
M12 N1N454 DIN2 GVSS 0 nch W=1.8U L=0.24U
M10 N1N508 DIN5 Q 0 nch W=1.8U L=0.24U
M14 GVSS DIN6 N1N508 0 nch W=1.8U L=0.24U
M11 GVSS DIN7 Q 0 nch W=0.9U L=0.24U
M7 Q DIN7 N1N452 VDD pch W=8.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi222s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N453 0 nch W=1U L=0.24U
M1 N1N441 DIN6 VDD VDD pch W=3.76U L=0.24U
M2 VDD DIN5 N1N441 VDD pch W=3.76U L=0.24U
M3 N1N443 DIN4 N1N441 VDD pch W=3.46U L=0.24U
M4 N1N441 DIN3 N1N443 VDD pch W=3.46U L=0.24U
M5 Q DIN1 N1N443 VDD pch W=3.2U L=0.24U
M6 N1N443 DIN2 Q VDD pch W=3.2U L=0.24U
M10 N1N453 DIN2 GVSS 0 nch W=1.1U L=0.24U
M8 Q DIN3 N1N517 0 nch W=1U L=0.24U
M11 N1N517 DIN4 GVSS 0 nch W=1.1U L=0.24U
M9 N1N455 DIN5 Q 0 nch W=1U L=0.24U
M12 GVSS DIN6 N1N455 0 nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi222s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N453 0 nch W=1.2U L=0.24U
M1 N1N441 DIN6 VDD VDD pch W=4.6U L=0.24U
M2 VDD DIN5 N1N441 VDD pch W=4.6U L=0.24U
M3 N1N443 DIN4 N1N441 VDD pch W=4.2U L=0.24U
M4 N1N441 DIN3 N1N443 VDD pch W=4.2U L=0.24U
M5 Q DIN1 N1N443 VDD pch W=3.8U L=0.24U
M6 N1N443 DIN2 Q VDD pch W=3.8U L=0.24U
M10 N1N453 DIN2 GVSS 0 nch W=1.4U L=0.24U
M8 Q DIN3 N1N474 0 nch W=1.2U L=0.24U
M11 N1N474 DIN4 GVSS 0 nch W=1.4U L=0.24U
M9 N1N455 DIN5 Q 0 nch W=1.2U L=0.24U
M12 GVSS DIN6 N1N455 0 nch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi222s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N449 DIN1 N1N453 0 nch W=1.3U L=0.24U
M1 N1N441 DIN6 VDD VDD pch W=3.8U L=0.24U
M3 N1N443 DIN4 N1N441 VDD pch W=3.6U L=0.24U
M5 N1N449 DIN1 N1N443 VDD pch W=3.3U L=0.24U
M2 VDD DIN5 N1N441 VDD pch W=3.8U L=0.24U
M4 N1N441 DIN3 N1N443 VDD pch W=3.6U L=0.24U
M6 N1N443 DIN2 N1N449 VDD pch W=3.3U L=0.24U
M10 N1N453 DIN2 GVSS 0 nch W=1.3U L=0.24U
M8 N1N449 DIN3 N1N474 0 nch W=1.3U L=0.24U
M11 N1N474 DIN4 GVSS 0 nch W=1.3U L=0.24U
M9 N1N455 DIN5 N1N449 0 nch W=1.3U L=0.24U
M12 GVSS DIN6 N1N455 0 nch W=1.3U L=0.24U
M14 N1N517 N1N449 GVSS 0 nch W=1.6U L=0.24U
M13 N1N517 N1N449 VDD VDD pch W=2.8U L=0.24U
M15 Q N1N517 VDD VDD pch W=4.7U L=0.24U
M16 Q N1N517 GVSS 0 nch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi22s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N445 0 nch W=1U L=0.24U
M1 N1N477 DIN3 VDD VDD pch W=2.6U L=0.24U
M3 Q DIN1 N1N477 VDD pch W=2.6U L=0.24U
M2 VDD DIN4 N1N477 VDD pch W=2.6U L=0.24U
M4 N1N477 DIN2 Q VDD pch W=2.6U L=0.24U
M7 N1N445 DIN2 GVSS 0 nch W=1U L=0.24U
M6 N1N447 DIN3 Q 0 nch W=1U L=0.24U
M8 GVSS DIN4 N1N447 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi22s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N445 0 nch W=1.3U L=0.24U
M1 N1N477 DIN3 VDD VDD pch W=3.3U L=0.24U
M3 Q DIN1 N1N477 VDD pch W=3.3U L=0.24U
M2 VDD DIN4 N1N477 VDD pch W=3.3U L=0.24U
M4 N1N477 DIN2 Q VDD pch W=3.3U L=0.24U
M7 N1N445 DIN2 GVSS 0 nch W=1.3U L=0.24U
M6 N1N447 DIN3 Q 0 nch W=1.3U L=0.24U
M8 GVSS DIN4 N1N447 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi22s3 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N445 0 nch W=1.84U L=0.24U
M1 N1N477 DIN3 VDD VDD pch W=4.6U L=0.24U
M3 Q DIN1 N1N477 VDD pch W=4.6U L=0.24U
M2 VDD DIN4 N1N477 VDD pch W=4.6U L=0.24U
M4 N1N477 DIN2 Q VDD pch W=4.6U L=0.24U
M7 N1N445 DIN2 GVSS 0 nch W=1.84U L=0.24U
M6 N1N447 DIN3 Q 0 nch W=1.84U L=0.24U
M8 GVSS DIN4 N1N447 0 nch W=1.84U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi23s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N497 0 nch W=1U L=0.24U
M1 N1N487 DIN3 VDD VDD pch W=2.66U L=0.24U
M3 VDD DIN5 N1N487 VDD pch W=2.66U L=0.24U
M5 N1N487 DIN2 Q VDD pch W=2.6U L=0.24U
M4 Q DIN1 N1N487 VDD pch W=2.6U L=0.24U
M7 N1N497 DIN2 GVSS 0 nch W=1U L=0.24U
M10 GVSS DIN5 N1N501 0 nch W=1.3U L=0.24U
M9 N1N501 DIN4 N1N499 0 nch W=1.3U L=0.24U
M8 N1N499 DIN3 Q 0 nch W=1.3U L=0.24U
M2 VDD DIN4 N1N487 VDD pch W=2.66U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi23s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M2 VDD DIN4 N1N435 VDD pch W=3.5U L=0.24U
M1 N1N435 DIN3 VDD VDD pch W=3.5U L=0.24U
M5 N1N435 DIN2 Q VDD pch W=3.4U L=0.24U
M4 Q DIN1 N1N435 VDD pch W=3.4U L=0.24U
M3 VDD DIN5 N1N435 VDD pch W=3.5U L=0.24U
M6 Q DIN1 N1N463 0 nch W=1.4U L=0.24U
M7 N1N463 DIN2 GVSS 0 nch W=1.4U L=0.24U
M10 GVSS DIN5 N1N467 0 nch W=1.8U L=0.24U
M8 N1N465 DIN3 Q 0 nch W=1.7U L=0.24U
M9 N1N467 DIN4 N1N465 0 nch W=1.76U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi23s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M2 VDD DIN4 N1N435 VDD pch W=4.8U L=0.24U
M1 N1N435 DIN3 VDD VDD pch W=4.8U L=0.24U
M5 N1N435 DIN2 Q VDD pch W=4.6U L=0.24U
M4 Q DIN1 N1N435 VDD pch W=4.6U L=0.24U
M3 VDD DIN5 N1N435 VDD pch W=4.8U L=0.24U
M6 Q DIN1 N1N463 0 nch W=1.9U L=0.24U
M7 N1N463 DIN2 GVSS 0 nch W=1.9U L=0.24U
M10 GVSS DIN5 N1N467 0 nch W=2.5U L=0.24U
M8 N1N465 DIN3 Q 0 nch W=2.3U L=0.24U
M9 N1N467 DIN4 N1N465 0 nch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi33s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN6 N1N481 0 nch W=1.7U L=0.24U
M1 N1N459 DIN2 VDD VDD pch W=2.56U L=0.24U
M4 Q DIN5 N1N459 VDD pch W=2.4U L=0.24U
M2 N1N459 DIN3 VDD VDD pch W=2.56U L=0.24U
M5 Q DIN6 N1N459 VDD pch W=2.4U L=0.24U
M3 VDD DIN1 N1N459 VDD pch W=2.56U L=0.24U
M6 N1N459 DIN4 Q VDD pch W=2.4U L=0.24U
M9 N1N481 DIN5 N1N483 0 nch W=1.7U L=0.24U
M11 N1N483 DIN4 GVSS 0 nch W=1.7U L=0.24U
M10 N1N487 DIN2 N1N485 0 nch W=1.7U L=0.24U
M8 Q DIN3 N1N485 0 nch W=1.7U L=0.24U
M12 GVSS DIN1 N1N487 0 nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi33s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN6 N1N481 0 nch W=2U L=0.24U
M1 N1N459 DIN2 VDD VDD pch W=3.5U L=0.24U
M2 N1N459 DIN3 VDD VDD pch W=3.5U L=0.24U
M4 Q DIN5 N1N459 VDD pch W=3.4U L=0.24U
M5 Q DIN6 N1N459 VDD pch W=3.4U L=0.24U
M3 VDD DIN1 N1N459 VDD pch W=3.5U L=0.24U
M6 N1N459 DIN4 Q VDD pch W=3.4U L=0.24U
M9 N1N481 DIN5 N1N483 0 nch W=2.5U L=0.24U
M11 N1N483 DIN4 GVSS 0 nch W=2.9U L=0.24U
M10 N1N487 DIN2 N1N485 0 nch W=2.5U L=0.24U
M8 Q DIN3 N1N485 0 nch W=2U L=0.24U
M12 GVSS DIN1 N1N487 0 nch W=2.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi33s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN6 N1N481 0 nch W=2.6U L=0.24U
M1 N1N459 DIN2 VDD VDD pch W=4.6U L=0.24U
M4 Q DIN5 N1N459 VDD pch W=4.4U L=0.24U
M2 N1N459 DIN3 VDD VDD pch W=4.6U L=0.24U
M5 Q DIN6 N1N459 VDD pch W=4.4U L=0.24U
M3 VDD DIN1 N1N459 VDD pch W=4.6U L=0.24U
M6 N1N459 DIN4 Q VDD pch W=4.4U L=0.24U
M8 Q DIN3 N1N485 0 nch W=2.6U L=0.24U
M11 N1N483 DIN4 GVSS 0 nch W=3.9U L=0.24U
M10 N1N487 DIN2 N1N485 0 nch W=3.4U L=0.24U
M9 N1N481 DIN5 N1N483 0 nch W=3.4U L=0.24U
M12 GVSS DIN1 N1N487 0 nch W=3.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi4111s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 Q DIN7 GVSS 0 nch W=0.6U L=0.24U
M5 N1N440 DIN7 N1N613 VDD pch W=5.4U L=0.24U
M6 N1N472 DIN6 N1N440 VDD pch W=5.2U L=0.24U
M7 Q DIN5 N1N472 VDD pch W=5U L=0.24U
M1 N1N613 DIN1 VDD VDD pch W=5.6U L=0.24U
M2 N1N613 DIN2 VDD VDD pch W=5.6U L=0.24U
M3 N1N613 DIN3 VDD VDD pch W=5.6U L=0.24U
M4 N1N613 DIN4 VDD VDD pch W=5.6U L=0.24U
M9 Q DIN6 GVSS 0 nch W=0.6U L=0.24U
M10 Q DIN5 GVSS 0 nch W=0.6U L=0.24U
M11 Q DIN4 N1N514 0 nch W=2.4U L=0.24U
M13 N1N515 DIN2 N1N501 0 nch W=2.4U L=0.24U
M14 N1N501 DIN1 GVSS 0 nch W=2.4U L=0.24U
M12 N1N515 DIN3 N1N514 0 nch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi4111s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 Q DIN7 GVSS 0 nch W=0.7U L=0.24U
M5 N1N440 DIN7 N1N613 VDD pch W=6.2U L=0.24U
M6 N1N472 DIN6 N1N440 VDD pch W=6U L=0.24U
M7 Q DIN5 N1N472 VDD pch W=5.8U L=0.24U
M1 N1N613 DIN1 VDD VDD pch W=6.3U L=0.24U
M2 N1N613 DIN2 VDD VDD pch W=6.3U L=0.24U
M3 N1N613 DIN3 VDD VDD pch W=6.3U L=0.24U
M4 N1N613 DIN4 VDD VDD pch W=6.3U L=0.24U
M9 Q DIN6 GVSS 0 nch W=0.7U L=0.24U
M10 Q DIN5 GVSS 0 nch W=0.7U L=0.24U
M11 Q DIN4 N1N514 0 nch W=2.8U L=0.24U
M13 N1N515 DIN2 N1N501 0 nch W=2.8U L=0.24U
M14 N1N501 DIN1 GVSS 0 nch W=2.8U L=0.24U
M12 N1N515 DIN3 N1N514 0 nch W=2.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi4111s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 N1N449 DIN7 GVSS 0 nch W=0.6U L=0.24U
M5 N1N440 DIN7 N1N639 VDD pch W=4.8U L=0.24U
M6 N1N472 DIN6 N1N440 VDD pch W=4.6U L=0.24U
M7 N1N449 DIN5 N1N472 VDD pch W=4.4U L=0.24U
M1 N1N639 DIN1 VDD VDD pch W=5U L=0.24U
M2 N1N639 DIN2 VDD VDD pch W=5U L=0.24U
M3 N1N639 DIN3 VDD VDD pch W=5U L=0.24U
M4 N1N639 DIN4 VDD VDD pch W=5U L=0.24U
M9 N1N449 DIN6 GVSS 0 nch W=0.6U L=0.24U
M10 N1N449 DIN5 GVSS 0 nch W=0.6U L=0.24U
M11 N1N449 DIN4 N1N514 0 nch W=2.4U L=0.24U
M13 N1N515 DIN2 N1N501 0 nch W=2.4U L=0.24U
M14 N1N501 DIN1 GVSS 0 nch W=2.4U L=0.24U
M12 N1N515 DIN3 N1N514 0 nch W=2.4U L=0.24U
M16 N1N591 N1N449 GVSS 0 nch W=2.2U L=0.24U
M15 N1N591 N1N449 VDD VDD pch W=4.8U L=0.24U
M17 Q N1N591 VDD VDD pch W=6.6U L=0.24U
M18 Q N1N591 GVSS 0 nch W=3.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi42s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N447 0 nch W=1.9U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=2.6U L=0.24U
M2 N1N440 DIN2 VDD VDD pch W=2.6U L=0.24U
M3 VDD DIN3 N1N440 VDD pch W=2.6U L=0.24U
M4 VDD DIN4 N1N440 VDD pch W=2.6U L=0.24U
M5 Q DIN5 N1N440 VDD pch W=2.6U L=0.24U
M6 N1N440 DIN6 Q VDD pch W=2.6U L=0.24U
M8 N1N447 DIN2 N1N463 0 nch W=1.9U L=0.24U
M9 N1N463 DIN3 N1N465 0 nch W=1.9U L=0.24U
M10 N1N465 DIN4 GVSS 0 nch W=1.9U L=0.24U
M11 N1N451 DIN5 Q 0 nch W=1U L=0.24U
M12 GVSS DIN6 N1N451 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi42s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N447 0 nch W=2.86U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=3.9U L=0.24U
M2 N1N440 DIN2 VDD VDD pch W=3.9U L=0.24U
M3 VDD DIN3 N1N440 VDD pch W=3.9U L=0.24U
M4 VDD DIN4 N1N440 VDD pch W=3.9U L=0.24U
M5 Q DIN5 N1N440 VDD pch W=3.9U L=0.24U
M6 N1N440 DIN6 Q VDD pch W=3.9U L=0.24U
M8 N1N447 DIN2 N1N463 0 nch W=2.86U L=0.24U
M9 N1N463 DIN3 N1N465 0 nch W=2.86U L=0.24U
M10 N1N465 DIN4 GVSS 0 nch W=2.86U L=0.24U
M11 N1N451 DIN5 Q 0 nch W=1.5U L=0.24U
M12 GVSS DIN6 N1N451 0 nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_aoi42s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N447 0 nch W=4.3U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=5.9U L=0.24U
M2 N1N440 DIN2 VDD VDD pch W=5.9U L=0.24U
M3 VDD DIN3 N1N440 VDD pch W=5.9U L=0.24U
M4 VDD DIN4 N1N440 VDD pch W=5.9U L=0.24U
M5 Q DIN5 N1N440 VDD pch W=5.9U L=0.24U
M6 N1N440 DIN6 Q VDD pch W=5.9U L=0.24U
M8 N1N447 DIN2 N1N463 0 nch W=4.3U L=0.24U
M9 N1N463 DIN3 N1N465 0 nch W=4.3U L=0.24U
M10 N1N465 DIN4 GVSS 0 nch W=4.3U L=0.24U
M11 N1N451 DIN5 Q 0 nch W=2.26U L=0.24U
M12 GVSS DIN6 N1N451 0 nch W=2.26U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_bshes1 INOUT1 INOUT2 E
M2 N1N313 E GVSS 0 nch W=0.8U L=0.24U
M1 N1N313 E VDD VDD pch W=1.2U L=0.24U
M3 INOUT2 N1N313 INOUT1 VDD pch W=1.2U L=0.24U
M4 INOUT1 E INOUT2 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_bshes2 INOUT2 E INOUT1
M2 N1N313 E GVSS 0 nch W=1U L=0.24U
M1 N1N313 E VDD VDD pch W=1.5U L=0.24U
M3 INOUT2 N1N313 INOUT1 VDD pch W=2.1U L=0.24U
M4 INOUT1 E INOUT2 0 nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_bshes3 INOUT2 E INOUT1
M2 N1N313 E GVSS 0 nch W=1.2U L=0.24U
M1 N1N313 E VDD VDD pch W=2U L=0.24U
M3 INOUT2 N1N313 INOUT1 VDD pch W=3.5U L=0.24U
M4 INOUT1 E INOUT2 0 nch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_bsles1 INOUT2 EB INOUT1
M2 N1N330 EB GVSS 0 nch W=0.9U L=0.24U
M1 N1N330 EB VDD VDD pch W=1.15U L=0.24U
M3 INOUT2 EB INOUT1 VDD pch W=1.45U L=0.24U
M4 INOUT1 N1N330 INOUT2 0 nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_bsles2 INOUT2 EB INOUT1
M2 N1N330 EB GVSS 0 nch W=1U L=0.24U
M1 N1N330 EB VDD VDD pch W=1.5U L=0.24U
M3 INOUT2 EB INOUT1 VDD pch W=2.1U L=0.24U
M4 INOUT1 N1N330 INOUT2 0 nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_bsles3 INOUT2 EB INOUT1
M2 N1N330 EB GVSS 0 nch W=1.2U L=0.24U
M1 N1N330 EB VDD VDD pch W=2U L=0.24U
M3 INOUT2 EB INOUT1 VDD pch W=3.5U L=0.24U
M4 INOUT1 N1N330 INOUT2 0 nch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_clc2s1 PIN0 CIN0 GIN0 GIN1 PIN1 OUTP OUTC OUTG
M14 OUTC N1N64 GVSS 0 nch W=0.72U L=0.24U
M7 OUTC N1N64 VDD VDD pch W=1.4U L=0.24U
M16 OUTG N1N145 GVSS 0 nch W=0.72U L=0.24U
M15 OUTG N1N145 VDD VDD pch W=1.4U L=0.24U
M17 N1N153 PIN0 VDD VDD pch W=0.9U L=0.24U
M18 N1N153 PIN1 VDD VDD pch W=0.9U L=0.24U
M19 N1N153 PIN0 N1N151 0 nch W=0.7U L=0.24U
M20 N1N151 PIN1 GVSS 0 nch W=0.7U L=0.24U
M22 OUTP N1N153 GVSS 0 nch W=0.9U L=0.24U
M21 OUTP N1N153 VDD VDD pch W=1.76U L=0.24U
M6 GVSS PIN0 N1N66 0 nch W=1.2U L=0.24U
M4 N1N64 GIN0 GVSS 0 nch W=0.6U L=0.24U
M5 N1N66 CIN0 N1N64 0 nch W=1.2U L=0.24U
M1 N1N60 PIN0 VDD VDD pch W=2.7U L=0.24U
M2 VDD CIN0 N1N60 VDD pch W=2.7U L=0.24U
M3 N1N64 GIN0 N1N60 VDD pch W=2.7U L=0.24U
M8 N1N86 GIN0 VDD VDD pch W=2.7U L=0.24U
M9 VDD PIN1 N1N86 VDD pch W=2.7U L=0.24U
M10 N1N145 GIN1 N1N86 VDD pch W=2.7U L=0.24U
M11 N1N145 GIN1 GVSS 0 nch W=0.6U L=0.24U
M12 N1N85 PIN1 N1N145 0 nch W=1.2U L=0.24U
M13 GVSS GIN0 N1N85 0 nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_clc2s2 PIN0 CIN0 GIN0 GIN1 PIN1 OUTP OUTC OUTG
M14 OUTC N1N64 GVSS 0 nch W=0.92U L=0.24U
M7 OUTC N1N64 VDD VDD pch W=1.7U L=0.24U
M16 OUTG N1N145 GVSS 0 nch W=0.92U L=0.24U
M15 OUTG N1N145 VDD VDD pch W=1.7U L=0.24U
M17 N1N153 PIN0 VDD VDD pch W=1.2U L=0.24U
M18 N1N153 PIN1 VDD VDD pch W=1.2U L=0.24U
M19 N1N153 PIN0 N1N151 0 nch W=0.9U L=0.24U
M20 N1N151 PIN1 GVSS 0 nch W=0.9U L=0.24U
M22 OUTP N1N153 GVSS 0 nch W=1.2U L=0.24U
M21 OUTP N1N153 VDD VDD pch W=2.26U L=0.24U
M6 GVSS PIN0 N1N66 0 nch W=1.6U L=0.24U
M4 N1N64 GIN0 GVSS 0 nch W=0.8U L=0.24U
M5 N1N66 CIN0 N1N64 0 nch W=1.6U L=0.24U
M1 N1N60 PIN0 VDD VDD pch W=3.5U L=0.24U
M2 VDD CIN0 N1N60 VDD pch W=3.5U L=0.24U
M3 N1N64 GIN0 N1N60 VDD pch W=3.5U L=0.24U
M8 N1N86 GIN0 VDD VDD pch W=3.5U L=0.24U
M9 VDD PIN1 N1N86 VDD pch W=3.5U L=0.24U
M10 N1N145 GIN1 N1N86 VDD pch W=3.5U L=0.24U
M11 N1N145 GIN1 GVSS 0 nch W=0.8U L=0.24U
M12 N1N85 PIN1 N1N145 0 nch W=1.6U L=0.24U
M13 GVSS GIN0 N1N85 0 nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_clc2s3 PIN0 CIN0 GIN0 GIN1 PIN1 OUTP OUTC OUTG
M14 OUTC N1N64 GVSS 0 nch W=1.26U L=0.24U
M7 OUTC N1N64 VDD VDD pch W=2.2U L=0.24U
M16 OUTG N1N145 GVSS 0 nch W=1.26U L=0.24U
M15 OUTG N1N145 VDD VDD pch W=2.2U L=0.24U
M17 N1N153 PIN0 VDD VDD pch W=1.74U L=0.24U
M18 N1N153 PIN1 VDD VDD pch W=1.74U L=0.24U
M19 N1N153 PIN0 N1N151 0 nch W=1.2U L=0.24U
M20 N1N151 PIN1 GVSS 0 nch W=1.2U L=0.24U
M22 OUTP N1N153 GVSS 0 nch W=1.5U L=0.24U
M21 OUTP N1N153 VDD VDD pch W=2.9U L=0.24U
M6 GVSS PIN0 N1N66 0 nch W=2U L=0.24U
M4 N1N64 GIN0 GVSS 0 nch W=1U L=0.24U
M5 N1N66 CIN0 N1N64 0 nch W=2U L=0.24U
M1 N1N60 PIN0 VDD VDD pch W=4.9U L=0.24U
M2 VDD CIN0 N1N60 VDD pch W=4.9U L=0.24U
M3 N1N64 GIN0 N1N60 VDD pch W=4.7U L=0.24U
M8 N1N86 GIN0 VDD VDD pch W=4.9U L=0.24U
M9 VDD PIN1 N1N86 VDD pch W=4.9U L=0.24U
M10 N1N145 GIN1 N1N86 VDD pch W=4.7U L=0.24U
M11 N1N145 GIN1 GVSS 0 nch W=1U L=0.24U
M12 N1N85 PIN1 N1N145 0 nch W=2U L=0.24U
M13 GVSS GIN0 N1N85 0 nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dchei24s1 BIN0 BIN1 E OUTD0 OUTD1 OUTD2 OUTD3
M15 OUTD1 N1N430 VDD VDD pch W=1.3U L=0.24U
M17 OUTD1 N1N301 VDD VDD pch W=1.3U L=0.24U
M20 N1N293 N1N301 GVSS 0 nch W=1.16U L=0.24U
M19 N1N294 BIN0 N1N293 0 nch W=1.16U L=0.24U
M18 OUTD1 N1N430 N1N294 0 nch W=1.16U L=0.24U
M16 OUTD1 BIN0 VDD VDD pch W=1.3U L=0.24U
M21 OUTD2 N1N430 VDD VDD pch W=1.3U L=0.24U
M23 OUTD2 BIN1 VDD VDD pch W=1.3U L=0.24U
M26 N1N325 BIN1 GVSS 0 nch W=1.16U L=0.24U
M25 N1N324 N1N290 N1N325 0 nch W=1.16U L=0.24U
M24 OUTD2 N1N430 N1N324 0 nch W=1.16U L=0.24U
M22 OUTD2 N1N290 VDD VDD pch W=1.3U L=0.24U
M9 OUTD0 N1N430 VDD VDD pch W=1.3U L=0.24U
M11 OUTD0 N1N301 VDD VDD pch W=1.3U L=0.24U
M14 N1N344 N1N301 GVSS 0 nch W=1.16U L=0.24U
M13 N1N343 N1N290 N1N344 0 nch W=1.16U L=0.24U
M12 OUTD0 N1N430 N1N343 0 nch W=1.16U L=0.24U
M10 OUTD0 N1N290 VDD VDD pch W=1.3U L=0.24U
M27 OUTD3 N1N430 VDD VDD pch W=1.3U L=0.24U
M29 OUTD3 BIN1 VDD VDD pch W=1.3U L=0.24U
M32 N1N363 BIN1 GVSS 0 nch W=1.16U L=0.24U
M31 N1N362 BIN0 N1N363 0 nch W=1.16U L=0.24U
M30 OUTD3 N1N430 N1N362 0 nch W=1.16U L=0.24U
M28 OUTD3 BIN0 VDD VDD pch W=1.3U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M2 N1N301 BIN1 GVSS 0 nch W=0.9U L=0.24U
M3 N1N290 BIN0 VDD VDD pch W=1.8U L=0.24U
M4 N1N290 BIN0 GVSS 0 nch W=0.9U L=0.24U
M5 N1N384 E VDD VDD pch W=1.2U L=0.24U
M7 N1N430 N1N384 VDD VDD pch W=1.6U L=0.24U
M6 N1N384 E GVSS 0 nch W=0.6U L=0.24U
M8 N1N430 N1N384 GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dchei24s2 BIN0 BIN1 E OUTD0 OUTD1 OUTD2 OUTD3
M15 OUTD1 N1N430 VDD VDD pch W=2U L=0.24U
M17 OUTD1 N1N301 VDD VDD pch W=2U L=0.24U
M20 N1N293 N1N301 GVSS 0 nch W=1.86U L=0.24U
M19 N1N294 BIN0 N1N293 0 nch W=1.86U L=0.24U
M18 OUTD1 N1N430 N1N294 0 nch W=1.86U L=0.24U
M16 OUTD1 BIN0 VDD VDD pch W=2U L=0.24U
M21 OUTD2 N1N430 VDD VDD pch W=2U L=0.24U
M23 OUTD2 BIN1 VDD VDD pch W=2U L=0.24U
M26 N1N325 BIN1 GVSS 0 nch W=1.86U L=0.24U
M25 N1N324 N1N290 N1N325 0 nch W=1.86U L=0.24U
M24 OUTD2 N1N430 N1N324 0 nch W=1.86U L=0.24U
M22 OUTD2 N1N290 VDD VDD pch W=2U L=0.24U
M9 OUTD0 N1N430 VDD VDD pch W=2U L=0.24U
M11 OUTD0 N1N301 VDD VDD pch W=2U L=0.24U
M14 N1N344 N1N301 GVSS 0 nch W=1.86U L=0.24U
M13 N1N343 N1N290 N1N344 0 nch W=1.86U L=0.24U
M12 OUTD0 N1N430 N1N343 0 nch W=1.86U L=0.24U
M10 OUTD0 N1N290 VDD VDD pch W=2U L=0.24U
M27 OUTD3 N1N430 VDD VDD pch W=2U L=0.24U
M29 OUTD3 BIN1 VDD VDD pch W=2U L=0.24U
M32 N1N363 BIN1 GVSS 0 nch W=1.86U L=0.24U
M31 N1N362 BIN0 N1N363 0 nch W=1.86U L=0.24U
M30 OUTD3 N1N430 N1N362 0 nch W=1.86U L=0.24U
M28 OUTD3 BIN0 VDD VDD pch W=2U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M2 N1N301 BIN1 GVSS 0 nch W=0.8U L=0.24U
M3 N1N290 BIN0 VDD VDD pch W=1.8U L=0.24U
M4 N1N290 BIN0 GVSS 0 nch W=0.9U L=0.24U
M5 N1N384 E VDD VDD pch W=1.2U L=0.24U
M7 N1N430 N1N384 VDD VDD pch W=1.6U L=0.24U
M6 N1N384 E GVSS 0 nch W=0.6U L=0.24U
M8 N1N430 N1N384 GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dchei24s3 BIN0 BIN1 E OUTD0 OUTD1 OUTD2 OUTD3
M15 OUTD1 N1N430 VDD VDD pch W=3U L=0.24U
M17 OUTD1 N1N301 VDD VDD pch W=3U L=0.24U
M20 N1N293 N1N301 GVSS 0 nch W=2.92U L=0.24U
M19 N1N294 BIN0 N1N293 0 nch W=2.92U L=0.24U
M18 OUTD1 N1N430 N1N294 0 nch W=2.92U L=0.24U
M16 OUTD1 BIN0 VDD VDD pch W=3U L=0.24U
M21 OUTD2 N1N430 VDD VDD pch W=3U L=0.24U
M23 OUTD2 BIN1 VDD VDD pch W=3U L=0.24U
M26 N1N325 BIN1 GVSS 0 nch W=2.92U L=0.24U
M25 N1N324 N1N290 N1N325 0 nch W=2.92U L=0.24U
M24 OUTD2 N1N430 N1N324 0 nch W=2.92U L=0.24U
M22 OUTD2 N1N290 VDD VDD pch W=3U L=0.24U
M9 OUTD0 N1N430 VDD VDD pch W=3U L=0.24U
M11 OUTD0 N1N301 VDD VDD pch W=3U L=0.24U
M14 N1N344 N1N301 GVSS 0 nch W=2.92U L=0.24U
M13 N1N343 N1N290 N1N344 0 nch W=2.92U L=0.24U
M12 OUTD0 N1N430 N1N343 0 nch W=2.92U L=0.24U
M10 OUTD0 N1N290 VDD VDD pch W=3U L=0.24U
M27 OUTD3 N1N430 VDD VDD pch W=3U L=0.24U
M29 OUTD3 BIN1 VDD VDD pch W=3U L=0.24U
M32 N1N363 BIN1 GVSS 0 nch W=2.92U L=0.24U
M31 N1N362 BIN0 N1N363 0 nch W=2.92U L=0.24U
M30 OUTD3 N1N430 N1N362 0 nch W=2.92U L=0.24U
M28 OUTD3 BIN0 VDD VDD pch W=3U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M2 N1N301 BIN1 GVSS 0 nch W=0.8U L=0.24U
M3 N1N290 BIN0 VDD VDD pch W=1.8U L=0.24U
M4 N1N290 BIN0 GVSS 0 nch W=0.9U L=0.24U
M5 N1N384 E VDD VDD pch W=1.2U L=0.24U
M7 N1N430 N1N384 VDD VDD pch W=1.6U L=0.24U
M6 N1N384 E GVSS 0 nch W=0.6U L=0.24U
M8 N1N430 N1N384 GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dci24s1 OUTD0 OUTD1 OUTD2 OUTD3 BIN1 BIN0
M2 N1N301 BIN1 GVSS 0 nch W=0.9U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N404 BIN0 GVSS 0 nch W=0.9U L=0.24U
M3 N1N404 BIN0 VDD VDD pch W=1.8U L=0.24U
M5 OUTD0 N1N404 VDD VDD pch W=1.66U L=0.24U
M6 VDD N1N301 OUTD0 VDD pch W=1.66U L=0.24U
M7 OUTD0 N1N404 N1N344 0 nch W=1.2U L=0.24U
M8 N1N344 N1N301 GVSS 0 nch W=1.2U L=0.24U
M12 N1N341 N1N301 GVSS 0 nch W=1.2U L=0.24U
M11 OUTD1 BIN0 N1N341 0 nch W=1.2U L=0.24U
M10 VDD N1N301 OUTD1 VDD pch W=1.66U L=0.24U
M9 OUTD1 BIN0 VDD VDD pch W=1.66U L=0.24U
M16 N1N338 N1N404 GVSS 0 nch W=1.2U L=0.24U
M15 OUTD2 BIN1 N1N338 0 nch W=1.2U L=0.24U
M14 VDD N1N404 OUTD2 VDD pch W=1.66U L=0.24U
M13 OUTD2 BIN1 VDD VDD pch W=1.66U L=0.24U
M20 N1N335 BIN1 GVSS 0 nch W=1.2U L=0.24U
M19 OUTD3 BIN0 N1N335 0 nch W=1.2U L=0.24U
M18 VDD BIN1 OUTD3 VDD pch W=1.66U L=0.24U
M17 OUTD3 BIN0 VDD VDD pch W=1.66U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dci24s2 OUTD0 OUTD1 OUTD2 OUTD3 BIN1 BIN0
M2 N1N301 BIN1 GVSS 0 nch W=0.9U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N404 BIN0 GVSS 0 nch W=0.9U L=0.24U
M3 N1N404 BIN0 VDD VDD pch W=1.8U L=0.24U
M5 OUTD0 N1N404 VDD VDD pch W=2.3U L=0.24U
M6 VDD N1N301 OUTD0 VDD pch W=2.3U L=0.24U
M7 OUTD0 N1N404 N1N344 0 nch W=1.8U L=0.24U
M8 N1N344 N1N301 GVSS 0 nch W=1.8U L=0.24U
M12 N1N341 N1N301 GVSS 0 nch W=1.8U L=0.24U
M11 OUTD1 BIN0 N1N341 0 nch W=1.8U L=0.24U
M10 VDD N1N301 OUTD1 VDD pch W=2.3U L=0.24U
M9 OUTD1 BIN0 VDD VDD pch W=2.3U L=0.24U
M16 N1N338 N1N404 GVSS 0 nch W=1.8U L=0.24U
M15 OUTD2 BIN1 N1N338 0 nch W=1.8U L=0.24U
M14 VDD N1N404 OUTD2 VDD pch W=2.3U L=0.24U
M13 OUTD2 BIN1 VDD VDD pch W=2.3U L=0.24U
M20 N1N335 BIN1 GVSS 0 nch W=1.8U L=0.24U
M19 OUTD3 BIN0 N1N335 0 nch W=1.8U L=0.24U
M18 VDD BIN1 OUTD3 VDD pch W=2.3U L=0.24U
M17 OUTD3 BIN0 VDD VDD pch W=2.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dci24s3 OUTD0 OUTD1 OUTD2 OUTD3 BIN1 BIN0
M2 N1N301 BIN1 GVSS 0 nch W=0.9U L=0.24U
M1 N1N301 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N404 BIN0 GVSS 0 nch W=0.9U L=0.24U
M3 N1N404 BIN0 VDD VDD pch W=1.8U L=0.24U
M5 OUTD0 N1N404 VDD VDD pch W=4.2U L=0.24U
M6 VDD N1N301 OUTD0 VDD pch W=4.2U L=0.24U
M7 OUTD0 N1N404 N1N344 0 nch W=4U L=0.24U
M8 N1N344 N1N301 GVSS 0 nch W=4U L=0.24U
M12 N1N341 N1N301 GVSS 0 nch W=4U L=0.24U
M11 OUTD1 BIN0 N1N341 0 nch W=4U L=0.24U
M10 VDD N1N301 OUTD1 VDD pch W=4.2U L=0.24U
M9 OUTD1 BIN0 VDD VDD pch W=4.2U L=0.24U
M16 N1N338 N1N404 GVSS 0 nch W=4U L=0.24U
M15 OUTD2 BIN1 N1N338 0 nch W=4U L=0.24U
M14 VDD N1N404 OUTD2 VDD pch W=4.2U L=0.24U
M13 OUTD2 BIN1 VDD VDD pch W=4.2U L=0.24U
M20 N1N335 BIN1 GVSS 0 nch W=4U L=0.24U
M19 OUTD3 BIN0 N1N335 0 nch W=4U L=0.24U
M18 VDD BIN1 OUTD3 VDD pch W=4.2U L=0.24U
M17 OUTD3 BIN0 VDD VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dclei24s1 BIN0 BIN1 EB OUTD0 OUTD1 OUTD2 OUTD3
M10 OUTD0 N1N344 N1N340 0 nch W=1.16U L=0.24U
M7 OUTD0 N1N344 VDD VDD pch W=1.3U L=0.24U
M8 OUTD0 N1N334 VDD VDD pch W=1.3U L=0.24U
M9 OUTD0 N1N346 VDD VDD pch W=1.3U L=0.24U
M11 N1N340 N1N334 N1N342 0 nch W=1.16U L=0.24U
M12 N1N342 N1N346 GVSS 0 nch W=1.16U L=0.24U
M16 OUTD1 N1N344 N1N373 0 nch W=1.16U L=0.24U
M13 OUTD1 N1N344 VDD VDD pch W=1.3U L=0.24U
M15 OUTD1 N1N346 VDD VDD pch W=1.3U L=0.24U
M14 OUTD1 BIN0 VDD VDD pch W=1.3U L=0.24U
M17 N1N373 BIN0 N1N374 0 nch W=1.16U L=0.24U
M18 N1N374 N1N346 GVSS 0 nch W=1.16U L=0.24U
M22 OUTD2 N1N344 N1N389 0 nch W=1.16U L=0.24U
M19 OUTD2 N1N344 VDD VDD pch W=1.3U L=0.24U
M21 OUTD2 BIN1 VDD VDD pch W=1.3U L=0.24U
M20 OUTD2 N1N334 VDD VDD pch W=1.3U L=0.24U
M23 N1N389 N1N334 N1N451 0 nch W=1.16U L=0.24U
M24 N1N451 BIN1 GVSS 0 nch W=1.16U L=0.24U
M28 OUTD3 N1N344 N1N405 0 nch W=1.16U L=0.24U
M25 OUTD3 N1N344 VDD VDD pch W=1.3U L=0.24U
M27 OUTD3 BIN1 VDD VDD pch W=1.3U L=0.24U
M26 OUTD3 BIN0 VDD VDD pch W=1.3U L=0.24U
M29 N1N405 BIN0 N1N406 0 nch W=1.16U L=0.24U
M30 N1N406 BIN1 GVSS 0 nch W=1.16U L=0.24U
M3 N1N346 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N346 BIN1 GVSS 0 nch W=0.9U L=0.24U
M1 N1N334 BIN0 VDD VDD pch W=1.8U L=0.24U
M2 N1N334 BIN0 GVSS 0 nch W=0.9U L=0.24U
M6 N1N344 EB GVSS 0 nch W=1.2U L=0.24U
M5 N1N344 EB VDD VDD pch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dclei24s2 BIN0 BIN1 EB OUTD0 OUTD1 OUTD2 OUTD3
M10 OUTD0 N1N344 N1N340 0 nch W=1.86U L=0.24U
M7 OUTD0 N1N344 VDD VDD pch W=2U L=0.24U
M8 OUTD0 N1N334 VDD VDD pch W=2U L=0.24U
M9 OUTD0 N1N346 VDD VDD pch W=2U L=0.24U
M11 N1N340 N1N334 N1N342 0 nch W=1.86U L=0.24U
M12 N1N342 N1N346 GVSS 0 nch W=1.86U L=0.24U
M16 OUTD1 N1N344 N1N373 0 nch W=1.86U L=0.24U
M13 OUTD1 N1N344 VDD VDD pch W=2U L=0.24U
M15 OUTD1 N1N346 VDD VDD pch W=2U L=0.24U
M14 OUTD1 BIN0 VDD VDD pch W=2U L=0.24U
M17 N1N373 BIN0 N1N374 0 nch W=1.86U L=0.24U
M18 N1N374 N1N346 GVSS 0 nch W=1.86U L=0.24U
M22 OUTD2 N1N344 N1N389 0 nch W=1.86U L=0.24U
M19 OUTD2 N1N344 VDD VDD pch W=2U L=0.24U
M21 OUTD2 BIN1 VDD VDD pch W=2U L=0.24U
M20 OUTD2 N1N334 VDD VDD pch W=2U L=0.24U
M23 N1N389 N1N334 N1N451 0 nch W=1.86U L=0.24U
M24 N1N451 BIN1 GVSS 0 nch W=1.86U L=0.24U
M28 OUTD3 N1N344 N1N405 0 nch W=1.86U L=0.24U
M25 OUTD3 N1N344 VDD VDD pch W=2U L=0.24U
M27 OUTD3 BIN1 VDD VDD pch W=2U L=0.24U
M26 OUTD3 BIN0 VDD VDD pch W=2U L=0.24U
M29 N1N405 BIN0 N1N406 0 nch W=1.86U L=0.24U
M30 N1N406 BIN1 GVSS 0 nch W=1.86U L=0.24U
M3 N1N346 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N346 BIN1 GVSS 0 nch W=0.9U L=0.24U
M1 N1N334 BIN0 VDD VDD pch W=1.8U L=0.24U
M2 N1N334 BIN0 GVSS 0 nch W=0.9U L=0.24U
M6 N1N344 EB GVSS 0 nch W=1.2U L=0.24U
M5 N1N344 EB VDD VDD pch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dclei24s3 BIN0 BIN1 EB OUTD0 OUTD1 OUTD2 OUTD3
M10 OUTD0 N1N344 N1N340 0 nch W=2.94U L=0.24U
M7 OUTD0 N1N344 VDD VDD pch W=3U L=0.24U
M8 OUTD0 N1N334 VDD VDD pch W=3U L=0.24U
M9 OUTD0 N1N346 VDD VDD pch W=3U L=0.24U
M11 N1N340 N1N334 N1N342 0 nch W=2.94U L=0.24U
M12 N1N342 N1N346 GVSS 0 nch W=2.94U L=0.24U
M16 OUTD1 N1N344 N1N373 0 nch W=2.94U L=0.24U
M13 OUTD1 N1N344 VDD VDD pch W=3U L=0.24U
M15 OUTD1 N1N346 VDD VDD pch W=3U L=0.24U
M14 OUTD1 BIN0 VDD VDD pch W=3U L=0.24U
M17 N1N373 BIN0 N1N374 0 nch W=2.94U L=0.24U
M18 N1N374 N1N346 GVSS 0 nch W=2.94U L=0.24U
M22 OUTD2 N1N344 N1N389 0 nch W=2.94U L=0.24U
M19 OUTD2 N1N344 VDD VDD pch W=3U L=0.24U
M21 OUTD2 BIN1 VDD VDD pch W=3U L=0.24U
M20 OUTD2 N1N334 VDD VDD pch W=3U L=0.24U
M23 N1N389 N1N334 N1N451 0 nch W=2.94U L=0.24U
M24 N1N451 BIN1 GVSS 0 nch W=2.94U L=0.24U
M28 OUTD3 N1N344 N1N405 0 nch W=2.94U L=0.24U
M25 OUTD3 N1N344 VDD VDD pch W=3U L=0.24U
M27 OUTD3 BIN1 VDD VDD pch W=3U L=0.24U
M26 OUTD3 BIN0 VDD VDD pch W=3U L=0.24U
M29 N1N405 BIN0 N1N406 0 nch W=2.94U L=0.24U
M30 N1N406 BIN1 GVSS 0 nch W=2.94U L=0.24U
M3 N1N346 BIN1 VDD VDD pch W=1.8U L=0.24U
M4 N1N346 BIN1 GVSS 0 nch W=0.9U L=0.24U
M1 N1N334 BIN0 VDD VDD pch W=1.8U L=0.24U
M2 N1N334 BIN0 GVSS 0 nch W=0.9U L=0.24U
M6 N1N344 EB GVSS 0 nch W=1.2U L=0.24U
M5 N1N344 EB VDD VDD pch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffacs1 Q QN CLRB CLK DIN
M17 TP7 CLRB VDD VDD pch W=1.3U L=0.24U
M21 Q TP8 VDD VDD pch W=3.14U L=0.24U
M9 TP5 TP3 VDD VDD pch W=1.3U L=0.24U
M24 QN Q GVSS 0 nch W=1.42U L=0.24U
M3 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M4 DIN TP1 TP3 0 nch W=0.8U L=0.24U
M13 TP5 CLK TP8 0 nch W=0.96U L=0.24U
M14 TP8 TP1 TP5 VDD pch W=1.4U L=0.24U
M6 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M15 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M16 TP8 TP1 TP7 0 nch W=0.8U L=0.24U
M23 QN Q VDD VDD pch W=3.02U L=0.24U
M5 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M11 TP5 TP3 TP6 0 nch W=0.9U L=0.24U
M19 TP7 Q TP9 0 nch W=0.9U L=0.24U
M22 Q TP8 GVSS 0 nch W=1.96U L=0.24U
M10 TP5 CLRB VDD VDD pch W=1.3U L=0.24U
M8 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M12 TP6 CLRB GVSS 0 nch W=0.9U L=0.24U
M1 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M7 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M18 TP7 Q VDD VDD pch W=1.3U L=0.24U
M20 TP9 CLRB GVSS 0 nch W=0.9U L=0.24U
M2 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffacs2 Q QN CLRB CLK DIN
M17 TP7 CLRB VDD VDD pch W=1.3U L=0.24U
M21 Q TP8 VDD VDD pch W=6.2U L=0.24U
M9 TP5 TP3 VDD VDD pch W=1.84U L=0.24U
M24 QN Q GVSS 0 nch W=2.68U L=0.24U
M3 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M4 DIN TP1 TP3 0 nch W=0.8U L=0.24U
M13 TP5 CLK TP8 0 nch W=1.52U L=0.24U
M14 TP8 TP1 TP5 VDD pch W=1.9U L=0.24U
M6 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M15 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M16 TP8 TP1 TP7 0 nch W=0.8U L=0.24U
M23 QN Q VDD VDD pch W=6.16U L=0.24U
M5 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M11 TP5 TP3 TP6 0 nch W=1.48U L=0.24U
M19 TP7 Q TP9 0 nch W=0.9U L=0.24U
M22 Q TP8 GVSS 0 nch W=3.98U L=0.24U
M10 TP5 CLRB VDD VDD pch W=1.84U L=0.24U
M8 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M12 TP6 CLRB GVSS 0 nch W=1.48U L=0.24U
M1 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M7 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M18 TP7 Q VDD VDD pch W=1.3U L=0.24U
M20 TP9 CLRB GVSS 0 nch W=0.9U L=0.24U
M2 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffascs1 SETB CLRB DIN CLK QN Q
M4 TP2 TP4 VDD VDD pch W=1.8U L=0.24U
M12 TP6 CLK GVSS 0 nch W=0.8U L=0.24U
M3 TP2 TP0 VDD VDD pch W=1.8U L=0.24U
M2 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M8 TP1 CLRB GVSS 0 nch W=0.8U L=0.24U
M7 TP1 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP1 VDD VDD pch W=2.2U L=0.24U
M10 TP4 TP1 GVSS 0 nch W=1.4U L=0.24U
M38 QN Q GVSS 0 nch W=1.44U L=0.24U
M30 TP14 Q VDD VDD pch W=1.3U L=0.24U
M33 Q TP13 VDD VDD pch W=3.18U L=0.24U
M23 TP11 TP8 TP12 0 nch W=2.2U L=0.24U
M13 TP8 CLK DIN VDD pch W=1.3U L=0.24U
M14 DIN TP6 TP8 0 nch W=0.8U L=0.24U
M25 TP11 CLK TP13 0 nch W=2.2U L=0.24U
M26 TP13 TP6 TP11 VDD pch W=2.5U L=0.24U
M15 TP8 CLK TP9 0 nch W=0.8U L=0.24U
M16 TP9 TP6 TP8 VDD pch W=1.3U L=0.24U
M27 TP14 CLK TP13 VDD pch W=1.3U L=0.24U
M28 TP13 TP6 TP14 0 nch W=0.8U L=0.24U
M17 TP9 TP2 VDD VDD pch W=1.3U L=0.24U
M21 TP11 TP8 VDD VDD pch W=2.4U L=0.24U
M22 TP11 TP4 VDD VDD pch W=2.4U L=0.24U
M29 TP14 TP4 VDD VDD pch W=1.3U L=0.24U
M37 QN Q VDD VDD pch W=3.18U L=0.24U
M31 TP14 Q TP15 0 nch W=0.8U L=0.24U
M20 TP10 TP11 GVSS 0 nch W=0.8U L=0.24U
M32 TP15 TP4 GVSS 0 nch W=0.8U L=0.24U
M24 TP12 TP4 GVSS 0 nch W=2.2U L=0.24U
M36 TP16 TP13 GVSS 0 nch W=2.64U L=0.24U
M34 Q TP2 VDD VDD pch W=3.18U L=0.24U
M35 Q TP2 TP16 0 nch W=2.64U L=0.24U
M18 TP9 TP11 VDD VDD pch W=1.3U L=0.24U
M19 TP9 TP2 TP10 0 nch W=0.8U L=0.24U
M11 TP6 CLK VDD VDD pch W=1.4U L=0.24U
M5 TP2 TP0 TP3 0 nch W=1.3U L=0.24U
M6 TP3 TP4 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffascs2 SETB CLRB DIN CLK QN Q
M4 TP2 TP4 VDD VDD pch W=2.82U L=0.24U
M12 TP6 CLK GVSS 0 nch W=0.8U L=0.24U
M3 TP2 TP0 VDD VDD pch W=2.82U L=0.24U
M2 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M8 TP1 CLRB GVSS 0 nch W=0.8U L=0.24U
M7 TP1 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP1 VDD VDD pch W=2.7U L=0.24U
M10 TP4 TP1 GVSS 0 nch W=2.2U L=0.24U
M38 QN Q GVSS 0 nch W=2.88U L=0.24U
M30 TP14 Q VDD VDD pch W=1.3U L=0.24U
M33 Q TP13 VDD VDD pch W=6.26U L=0.24U
M23 TP11 TP8 TP12 0 nch W=2.92U L=0.24U
M13 TP8 CLK DIN VDD pch W=1.3U L=0.24U
M14 DIN TP6 TP8 0 nch W=0.8U L=0.24U
M25 TP11 CLK TP13 0 nch W=2.7U L=0.24U
M26 TP13 TP6 TP11 VDD pch W=3U L=0.24U
M15 TP8 CLK TP9 0 nch W=0.8U L=0.24U
M16 TP9 TP6 TP8 VDD pch W=1.3U L=0.24U
M27 TP14 CLK TP13 VDD pch W=1.3U L=0.24U
M28 TP13 TP6 TP14 0 nch W=0.8U L=0.24U
M17 TP9 TP2 VDD VDD pch W=1.3U L=0.24U
M21 TP11 TP8 VDD VDD pch W=3.24U L=0.24U
M22 TP11 TP4 VDD VDD pch W=3.24U L=0.24U
M29 TP14 TP4 VDD VDD pch W=1.3U L=0.24U
M37 QN Q VDD VDD pch W=6.2U L=0.24U
M31 TP14 Q TP15 0 nch W=0.8U L=0.24U
M20 TP10 TP11 GVSS 0 nch W=0.8U L=0.24U
M32 TP15 TP4 GVSS 0 nch W=0.8U L=0.24U
M24 TP12 TP4 GVSS 0 nch W=2.92U L=0.24U
M36 TP16 TP13 GVSS 0 nch W=5.26U L=0.24U
M34 Q TP2 VDD VDD pch W=6.26U L=0.24U
M35 Q TP2 TP16 0 nch W=5.26U L=0.24U
M18 TP9 TP11 VDD VDD pch W=1.3U L=0.24U
M19 TP9 TP2 TP10 0 nch W=0.8U L=0.24U
M11 TP6 CLK VDD VDD pch W=1.6U L=0.24U
M5 TP2 TP0 TP3 0 nch W=2.2U L=0.24U
M6 TP3 TP4 GVSS 0 nch W=2.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffass1 Q QN SETB CLK DIN
M19 TP7 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 DIN GVSS 0 nch W=0.8U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.3U L=0.24U
M23 QN TP8 VDD VDD pch W=3.14U L=0.24U
M11 TP5 TP3 VDD VDD pch W=1.3U L=0.24U
M26 Q QN GVSS 0 nch W=1.42U L=0.24U
M5 TP3 CLK TP0 VDD pch W=1.3U L=0.24U
M6 TP0 TP1 TP3 0 nch W=0.8U L=0.24U
M15 TP5 CLK TP8 0 nch W=0.96U L=0.24U
M16 TP8 TP1 TP5 VDD pch W=1.4U L=0.24U
M8 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M17 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M18 TP8 TP1 TP7 0 nch W=0.8U L=0.24U
M25 Q QN VDD VDD pch W=3.02U L=0.24U
M7 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M13 TP5 TP3 TP6 0 nch W=0.9U L=0.24U
M21 TP7 QN TP9 0 nch W=0.9U L=0.24U
M24 QN TP8 GVSS 0 nch W=1.96U L=0.24U
M12 TP5 SETB VDD VDD pch W=1.3U L=0.24U
M10 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M14 TP6 SETB GVSS 0 nch W=0.9U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M20 TP7 QN VDD VDD pch W=1.3U L=0.24U
M22 TP9 SETB GVSS 0 nch W=0.9U L=0.24U
M4 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffass2 Q QN SETB CLK DIN
M19 TP7 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 DIN GVSS 0 nch W=0.8U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.3U L=0.24U
M23 QN TP8 VDD VDD pch W=6.2U L=0.24U
M11 TP5 TP3 VDD VDD pch W=1.84U L=0.24U
M26 Q QN GVSS 0 nch W=2.68U L=0.24U
M5 TP3 CLK TP0 VDD pch W=1.3U L=0.24U
M6 TP0 TP1 TP3 0 nch W=0.8U L=0.24U
M15 TP5 CLK TP8 0 nch W=1.52U L=0.24U
M16 TP8 TP1 TP5 VDD pch W=1.9U L=0.24U
M8 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M17 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M18 TP8 TP1 TP7 0 nch W=0.8U L=0.24U
M25 Q QN VDD VDD pch W=6.16U L=0.24U
M7 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M13 TP5 TP3 TP6 0 nch W=1.48U L=0.24U
M21 TP7 QN TP9 0 nch W=0.9U L=0.24U
M24 QN TP8 GVSS 0 nch W=3.98U L=0.24U
M12 TP5 SETB VDD VDD pch W=1.84U L=0.24U
M10 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M14 TP6 SETB GVSS 0 nch W=1.48U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M20 TP7 QN VDD VDD pch W=1.3U L=0.24U
M22 TP9 SETB GVSS 0 nch W=0.9U L=0.24U
M4 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffcs1 Q QN CLK DIN CLRB
M8 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M9 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M10 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M15 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M17 TP6 CLK TP7 0 nch W=0.8U L=0.24U
M18 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M23 QN TP7 VDD VDD pch W=3.14U L=0.24U
M24 QN TP7 GVSS 0 nch W=2.06U L=0.24U
M11 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M12 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M14 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M19 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M25 Q QN VDD VDD pch W=2.94U L=0.24U
M26 Q QN GVSS 0 nch W=1.28U L=0.24U
M16 TP6 TP4 GVSS 0 nch W=0.8U L=0.24U
M7 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M22 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M20 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M21 TP8 QN VDD VDD pch W=1.3U L=0.24U
M3 TP2 DIN TP1 0 nch W=0.8U L=0.24U
M13 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M4 TP1 CLRB GVSS 0 nch W=0.8U L=0.24U
M2 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M1 TP2 DIN VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffcs2 Q QN CLK DIN CLRB
M8 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M9 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M10 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M15 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M17 TP6 CLK TP7 0 nch W=1.3U L=0.24U
M18 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M23 QN TP7 VDD VDD pch W=6.24U L=0.24U
M24 QN TP7 GVSS 0 nch W=3.98U L=0.24U
M11 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M12 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M14 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M19 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M25 Q QN VDD VDD pch W=5.92U L=0.24U
M26 Q QN GVSS 0 nch W=2.66U L=0.24U
M16 TP6 TP4 GVSS 0 nch W=1.26U L=0.24U
M7 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M22 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M20 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M21 TP8 QN VDD VDD pch W=1.3U L=0.24U
M3 TP2 DIN TP1 0 nch W=0.8U L=0.24U
M13 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M4 TP1 CLRB GVSS 0 nch W=0.8U L=0.24U
M2 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M1 TP2 DIN VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffles1 EB DIN CLK QN Q
M8 N1N80 TP7 GVSS 0 nch W=0.8U L=0.24U
M7 N1N80 TP7 VDD VDD pch W=1.3U L=0.24U
M12 TP21 TP1 TP3 0 nch W=0.8U L=0.24U
M19 TP5 CLK TP6 0 nch W=0.8U L=0.24U
M20 TP6 TP1 TP5 VDD pch W=1.3U L=0.24U
M26 Q TP6 GVSS 0 nch W=2.06U L=0.24U
M13 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M14 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M15 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M16 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M21 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M22 TP6 TP1 TP7 0 nch W=0.8U L=0.24U
M24 TP7 Q GVSS 0 nch W=0.8U L=0.24U
M28 QN Q GVSS 0 nch W=1.28U L=0.24U
M18 TP5 TP3 GVSS 0 nch W=0.8U L=0.24U
M11 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M17 TP5 TP3 VDD VDD pch W=1.8U L=0.24U
M27 QN Q VDD VDD pch W=2.94U L=0.24U
M25 Q TP6 VDD VDD pch W=3.14U L=0.24U
M9 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M23 TP7 Q VDD VDD pch W=1.3U L=0.24U
M10 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M3 N1N80 EB TP21 0 nch W=0.8U L=0.24U
M4 TP21 TP20 N1N80 VDD pch W=1.3U L=0.24U
M5 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M6 TP21 EB DIN VDD pch W=1.3U L=0.24U
M1 TP20 EB VDD VDD pch W=1.3U L=0.24U
M2 TP20 EB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffles2 EB DIN CLK QN Q
M8 N1N80 TP7 GVSS 0 nch W=0.8U L=0.24U
M7 N1N80 TP7 VDD VDD pch W=1.3U L=0.24U
M12 TP21 TP1 TP3 0 nch W=0.8U L=0.24U
M19 TP5 CLK TP6 0 nch W=1.3U L=0.24U
M20 TP6 TP1 TP5 VDD pch W=1.8U L=0.24U
M26 Q TP6 GVSS 0 nch W=3.98U L=0.24U
M13 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M14 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M15 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M16 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M21 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M22 TP6 TP1 TP7 0 nch W=0.8U L=0.24U
M24 TP7 Q GVSS 0 nch W=0.8U L=0.24U
M28 QN Q GVSS 0 nch W=2.66U L=0.24U
M18 TP5 TP3 GVSS 0 nch W=1.26U L=0.24U
M11 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M17 TP5 TP3 VDD VDD pch W=2.78U L=0.24U
M27 QN Q VDD VDD pch W=5.92U L=0.24U
M25 Q TP6 VDD VDD pch W=6.24U L=0.24U
M9 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M23 TP7 Q VDD VDD pch W=1.3U L=0.24U
M10 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M3 N1N80 EB TP21 0 nch W=0.8U L=0.24U
M4 TP21 TP20 N1N80 VDD pch W=1.3U L=0.24U
M5 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M6 TP21 EB DIN VDD pch W=1.3U L=0.24U
M1 TP20 EB VDD VDD pch W=1.3U L=0.24U
M2 TP20 EB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffs1 Q QN CLK DIN
M8 DIN TP1 TP3 0 nch W=0.8U L=0.24U
M15 TP5 CLK TP6 0 nch W=0.8U L=0.24U
M16 TP6 TP1 TP5 VDD pch W=1.3U L=0.24U
M20 Q TP6 GVSS 0 nch W=2.06U L=0.24U
M9 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M10 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M14 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M17 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M18 TP6 TP1 TP7 0 nch W=0.8U L=0.24U
M21 TP7 Q VDD VDD pch W=1.3U L=0.24U
M22 TP7 Q GVSS 0 nch W=0.8U L=0.24U
M24 QN Q GVSS 0 nch W=1.28U L=0.24U
M12 TP5 TP3 GVSS 0 nch W=0.8U L=0.24U
M7 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M11 TP5 TP3 VDD VDD pch W=1.8U L=0.24U
M23 QN Q VDD VDD pch W=2.94U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M19 Q TP6 VDD VDD pch W=3.14U L=0.24U
M4 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffs2 DIN CLK Q QN
M8 DIN TP1 TP3 0 nch W=0.8U L=0.24U
M15 TP5 CLK TP6 0 nch W=1.3U L=0.24U
M16 TP6 TP1 TP5 VDD pch W=1.8U L=0.24U
M20 Q TP6 GVSS 0 nch W=3.98U L=0.24U
M9 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M10 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M14 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M17 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M18 TP6 TP1 TP7 0 nch W=0.8U L=0.24U
M21 TP7 Q VDD VDD pch W=1.3U L=0.24U
M22 TP7 Q GVSS 0 nch W=0.8U L=0.24U
M24 QN Q GVSS 0 nch W=2.66U L=0.24U
M12 TP5 TP3 GVSS 0 nch W=1.26U L=0.24U
M7 TP3 CLK DIN VDD pch W=1.3U L=0.24U
M11 TP5 TP3 VDD VDD pch W=2.76U L=0.24U
M23 QN Q VDD VDD pch W=5.92U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M19 Q TP6 VDD VDD pch W=6.24U L=0.24U
M4 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffscs1 DIN SETB CLRB CLK Q OUTB
M11 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M12 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M17 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M19 TP6 CLK TP7 0 nch W=0.8U L=0.24U
M20 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M25 QN TP7 VDD VDD pch W=3.14U L=0.24U
M26 QN TP7 GVSS 0 nch W=2.06U L=0.24U
M13 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M14 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M16 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M21 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M27 Q QN VDD VDD pch W=2.94U L=0.24U
M28 Q QN GVSS 0 nch W=1.28U L=0.24U
M18 TP6 TP4 GVSS 0 nch W=0.8U L=0.24U
M9 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M10 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M24 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M22 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M23 TP8 QN VDD VDD pch W=1.3U L=0.24U
M15 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M4 TP2 DIN TP1 VDD pch W=1.3U L=0.24U
M5 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M6 TP2 CLRB TP9 0 nch W=0.8U L=0.24U
M7 TP9 DIN GVSS 0 nch W=0.8U L=0.24U
M8 TP9 TP0 GVSS 0 nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffscs2 DIN SETB CLRB CLK Q OUTB
M11 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M12 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M17 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M19 TP6 CLK TP7 0 nch W=1.3U L=0.24U
M20 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M25 QN TP7 VDD VDD pch W=6.24U L=0.24U
M26 QN TP7 GVSS 0 nch W=3.98U L=0.24U
M13 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M14 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M16 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M21 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M27 Q QN VDD VDD pch W=5.92U L=0.24U
M28 Q QN GVSS 0 nch W=2.66U L=0.24U
M18 TP6 TP4 GVSS 0 nch W=1.26U L=0.24U
M9 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M10 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M24 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M22 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M23 TP8 QN VDD VDD pch W=1.3U L=0.24U
M15 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M4 TP2 DIN TP1 VDD pch W=1.3U L=0.24U
M5 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M6 TP2 CLRB TP9 0 nch W=0.8U L=0.24U
M7 TP9 DIN GVSS 0 nch W=0.8U L=0.24U
M8 TP9 TP0 GVSS 0 nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffss1 SETB DIN CLK QN Q
M5 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M1 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M8 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M9 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M10 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M15 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M17 TP6 CLK TP7 0 nch W=0.8U L=0.24U
M18 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M23 QN TP7 VDD VDD pch W=3.14U L=0.24U
M24 QN TP7 GVSS 0 nch W=2.06U L=0.24U
M11 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M12 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M14 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M19 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M25 Q QN VDD VDD pch W=2.94U L=0.24U
M26 Q QN GVSS 0 nch W=1.28U L=0.24U
M16 TP6 TP4 GVSS 0 nch W=0.8U L=0.24U
M7 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M22 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M2 TP2 DIN TP1 VDD pch W=1.3U L=0.24U
M3 TP2 DIN GVSS 0 nch W=0.8U L=0.24U
M4 TP2 TP0 GVSS 0 nch W=0.8U L=0.24U
M20 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M21 TP8 QN VDD VDD pch W=1.3U L=0.24U
M13 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M6 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dffss2 SETB DIN CLK QN Q
M5 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M1 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M8 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M9 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M10 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M15 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M17 TP6 CLK TP7 0 nch W=1.3U L=0.24U
M18 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M23 QN TP7 VDD VDD pch W=6.24U L=0.24U
M24 QN TP7 GVSS 0 nch W=3.98U L=0.24U
M11 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M12 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M14 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M19 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M25 Q QN VDD VDD pch W=5.92U L=0.24U
M26 Q QN GVSS 0 nch W=2.66U L=0.24U
M16 TP6 TP4 GVSS 0 nch W=1.26U L=0.24U
M7 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M22 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M2 TP2 DIN TP1 VDD pch W=1.3U L=0.24U
M3 TP2 DIN GVSS 0 nch W=0.8U L=0.24U
M4 TP2 TP0 GVSS 0 nch W=0.8U L=0.24U
M20 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M21 TP8 QN VDD VDD pch W=1.3U L=0.24U
M13 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M6 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s1 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=1.8U L=0.24U
M4 GVSS DIN2 Q2 0 nch W=0.74U L=0.24U
M2 Q1 DIN1 GVSS 0 nch W=0.74U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s10 DIN1 DIN2 Q1 Q2
M1 N1N255 DIN1 VDD VDD pch W=9.5U L=0.24U
M2 N1N255 DIN1 GVSS 0 nch W=6.8U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=20.28U L=0.24U
M4 N1N266 N1N255 GVSS 0 nch W=14.56U L=0.24U
M5 Q1 N1N266 VDD VDD pch W=47.64U L=0.24U
M6 Q1 N1N266 GVSS 0 nch W=19.5U L=0.24U
M8 N1N340 DIN2 GVSS 0 nch W=6.8U L=0.24U
M7 N1N340 DIN2 VDD VDD pch W=9.5U L=0.24U
M10 N1N347 N1N340 GVSS 0 nch W=14.56U L=0.24U
M9 N1N347 N1N340 VDD VDD pch W=20.28U L=0.24U
M12 Q2 N1N347 GVSS 0 nch W=19.5U L=0.24U
M11 Q2 N1N347 VDD VDD pch W=47.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s11 DIN1 DIN2 Q1 Q2
M3 N1N255 N1N253 VDD VDD pch W=9U L=0.24U
M4 N1N255 N1N253 GVSS 0 nch W=4.5U L=0.24U
M5 N1N266 N1N255 VDD VDD pch W=20U L=0.24U
M6 N1N266 N1N255 GVSS 0 nch W=11U L=0.24U
M7 N1N268 N1N266 VDD VDD pch W=40U L=0.24U
M8 N1N268 N1N266 GVSS 0 nch W=26U L=0.24U
M1 N1N253 DIN1 VDD VDD pch W=4U L=0.24U
M2 N1N253 DIN1 GVSS 0 nch W=2.2U L=0.24U
M9 Q1 N1N268 VDD VDD pch W=84U L=0.24U
M10 Q1 N1N268 GVSS 0 nch W=42U L=0.24U
M14 N1N312 N1N299 GVSS 0 nch W=4.5U L=0.24U
M13 N1N312 N1N299 VDD VDD pch W=9U L=0.24U
M16 N1N319 N1N312 GVSS 0 nch W=11U L=0.24U
M15 N1N319 N1N312 VDD VDD pch W=20U L=0.24U
M18 N1N297 N1N319 GVSS 0 nch W=26U L=0.24U
M17 N1N297 N1N319 VDD VDD pch W=40U L=0.24U
M12 N1N299 DIN2 GVSS 0 nch W=2.2U L=0.24U
M11 N1N299 DIN2 VDD VDD pch W=4U L=0.24U
M20 Q2 N1N297 GVSS 0 nch W=42U L=0.24U
M19 Q2 N1N297 VDD VDD pch W=84U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s12 DIN1 DIN2 Q1 Q2
M3 N1N255 N1N253 VDD VDD pch W=16.5U L=0.24U
M4 N1N255 N1N253 GVSS 0 nch W=9.8U L=0.24U
M5 N1N266 N1N255 VDD VDD pch W=36.4U L=0.24U
M6 N1N266 N1N255 GVSS 0 nch W=20.6U L=0.24U
M7 N1N268 N1N266 VDD VDD pch W=88.3U L=0.24U
M8 N1N268 N1N266 GVSS 0 nch W=50.9U L=0.24U
M1 N1N253 DIN1 VDD VDD pch W=8.3U L=0.24U
M2 N1N253 DIN1 GVSS 0 nch W=5U L=0.24U
M9 Q1 N1N268 VDD VDD pch W=180.8U L=0.24U
M10 Q1 N1N268 GVSS 0 nch W=78.6U L=0.24U
M14 N1N312 N1N299 GVSS 0 nch W=9.8U L=0.24U
M13 N1N312 N1N299 VDD VDD pch W=16.5U L=0.24U
M16 N1N319 N1N312 GVSS 0 nch W=20.6U L=0.24U
M15 N1N319 N1N312 VDD VDD pch W=36.4U L=0.24U
M18 N1N297 N1N319 GVSS 0 nch W=50.9U L=0.24U
M17 N1N297 N1N319 VDD VDD pch W=88.3U L=0.24U
M12 N1N299 DIN2 GVSS 0 nch W=5U L=0.24U
M11 N1N299 DIN2 VDD VDD pch W=8.3U L=0.24U
M20 Q2 N1N297 GVSS 0 nch W=78.6U L=0.24U
M19 Q2 N1N297 VDD VDD pch W=180.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s2 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=3.16U L=0.24U
M4 GVSS DIN2 Q2 0 nch W=1.24U L=0.24U
M2 Q1 DIN1 GVSS 0 nch W=1.24U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=3.16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s3 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=4.98U L=0.24U
M4 GVSS DIN2 Q2 0 nch W=2.14U L=0.24U
M2 Q1 DIN1 GVSS 0 nch W=2.14U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=4.98U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s4 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=5.8U L=0.24U
M4 GVSS DIN2 Q2 0 nch W=2.5U L=0.24U
M2 Q1 DIN1 GVSS 0 nch W=2.5U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=5.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s5 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=8.28U L=0.24U
M4 GVSS DIN2 Q2 0 nch W=3.5U L=0.24U
M2 Q1 DIN1 GVSS 0 nch W=3.5U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=8.28U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s6 Q1 Q2 DIN1 DIN2
M3 VDD DIN2 Q2 VDD pch W=10.7U L=0.24U
M4 GVSS DIN2 Q2 0 nch W=4.7U L=0.24U
M2 Q1 DIN1 GVSS 0 nch W=4.7U L=0.24U
M1 Q1 DIN1 VDD VDD pch W=10.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s7 DIN1 DIN2 Q1 Q2
M1 N1N255 DIN1 VDD VDD pch W=4.1U L=0.24U
M2 N1N255 DIN1 GVSS 0 nch W=1.9U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=5.5U L=0.24U
M4 N1N266 N1N255 GVSS 0 nch W=3.1U L=0.24U
M5 Q1 N1N266 VDD VDD pch W=15.2U L=0.24U
M6 Q1 N1N266 GVSS 0 nch W=8.5U L=0.24U
M8 N1N340 DIN2 GVSS 0 nch W=1.9U L=0.24U
M7 N1N340 DIN2 VDD VDD pch W=4.1U L=0.24U
M10 N1N347 N1N340 GVSS 0 nch W=3.1U L=0.24U
M9 N1N347 N1N340 VDD VDD pch W=5.5U L=0.24U
M12 Q2 N1N347 GVSS 0 nch W=8.5U L=0.24U
M11 Q2 N1N347 VDD VDD pch W=15.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s8 DIN1 DIN2 Q1 Q2
M1 N1N255 DIN1 VDD VDD pch W=5.6U L=0.24U
M2 N1N255 DIN1 GVSS 0 nch W=4U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=12U L=0.24U
M4 N1N266 N1N255 GVSS 0 nch W=8.6U L=0.24U
M5 Q1 N1N266 VDD VDD pch W=25.4U L=0.24U
M6 Q1 N1N266 GVSS 0 nch W=12.7U L=0.24U
M8 N1N340 DIN2 GVSS 0 nch W=4U L=0.24U
M7 N1N340 DIN2 VDD VDD pch W=5.6U L=0.24U
M10 N1N347 N1N340 GVSS 0 nch W=8.6U L=0.24U
M9 N1N347 N1N340 VDD VDD pch W=12U L=0.24U
M12 Q2 N1N347 GVSS 0 nch W=12.7U L=0.24U
M11 Q2 N1N347 VDD VDD pch W=25.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_di2s9 DIN1 DIN2 Q1 Q2
M1 N1N255 DIN1 VDD VDD pch W=7.3U L=0.24U
M2 N1N255 DIN1 GVSS 0 nch W=5.2U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=15.6U L=0.24U
M4 N1N266 N1N255 GVSS 0 nch W=11.2U L=0.24U
M5 Q1 N1N266 VDD VDD pch W=35.8U L=0.24U
M6 Q1 N1N266 GVSS 0 nch W=15U L=0.24U
M8 N1N340 DIN2 GVSS 0 nch W=5.2U L=0.24U
M7 N1N340 DIN2 VDD VDD pch W=7.3U L=0.24U
M10 N1N347 N1N340 GVSS 0 nch W=11.2U L=0.24U
M9 N1N347 N1N340 VDD VDD pch W=15.6U L=0.24U
M12 Q2 N1N347 GVSS 0 nch W=15U L=0.24U
M11 Q2 N1N347 VDD VDD pch W=35.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dsmxc31s1 Q DIN1 CLK DIN2
M7 N1N280 DIN1 N1N270 0 nch W=0.6U L=0.24U
M3 N1N261 DIN2 VDD VDD pch W=1.1U L=0.24U
M5 N1N280 N1N276 N1N261 VDD pch W=1.1U L=0.24U
M4 VDD CLK N1N263 VDD pch W=1.1U L=0.24U
M6 N1N263 DIN1 N1N280 VDD pch W=1.1U L=0.24U
M9 N1N270 N1N276 GVSS 0 nch W=0.6U L=0.24U
M2 N1N276 CLK GVSS 0 nch W=0.6U L=0.24U
M1 N1N276 CLK VDD VDD pch W=1.2U L=0.24U
M8 N1N272 CLK N1N280 0 nch W=0.6U L=0.24U
M10 GVSS DIN2 N1N272 0 nch W=0.6U L=0.24U
M11 Q N1N280 VDD VDD pch W=1.84U L=0.24U
M12 Q N1N280 GVSS 0 nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_dsmxc31s2 Q DIN1 CLK DIN2
M7 N1N280 DIN1 N1N270 0 nch W=0.8U L=0.24U
M3 N1N261 DIN2 VDD VDD pch W=1.5U L=0.24U
M5 N1N280 N1N276 N1N261 VDD pch W=1.5U L=0.24U
M4 VDD CLK N1N263 VDD pch W=1.5U L=0.24U
M6 N1N263 DIN1 N1N280 VDD pch W=1.5U L=0.24U
M9 N1N270 N1N276 GVSS 0 nch W=0.8U L=0.24U
M2 N1N276 CLK GVSS 0 nch W=0.6U L=0.24U
M1 N1N276 CLK VDD VDD pch W=1.2U L=0.24U
M8 N1N272 CLK N1N280 0 nch W=0.8U L=0.24U
M10 GVSS DIN2 N1N272 0 nch W=0.8U L=0.24U
M11 Q N1N280 VDD VDD pch W=2.6U L=0.24U
M12 Q N1N280 GVSS 0 nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_fadd1s1 OUTS OUTC AIN BIN CIN
M1 TP9 AIN VDD VDD pch W=1.2U L=0.24U
M2 TP0 BIN TP9 VDD pch W=1.1U L=0.24U
M3 TP0 BIN TP8 0 nch W=0.8U L=0.24U
M4 TP8 AIN GVSS 0 nch W=0.9U L=0.24U
M5 TP10 AIN VDD VDD pch W=1.2U L=0.24U
M6 VDD BIN TP10 VDD pch W=1.2U L=0.24U
M7 TP10 CIN TP0 VDD pch W=1.1U L=0.24U
M8 TP11 CIN TP0 0 nch W=0.8U L=0.24U
M9 GVSS BIN TP11 0 nch W=0.9U L=0.24U
M10 TP11 AIN GVSS 0 nch W=0.9U L=0.24U
M11 TP1 AIN VDD VDD pch W=1.4U L=0.24U
M12 TP3 TP0 TP1 VDD pch W=1.1U L=0.24U
M13 TP3 TP0 TP2 0 nch W=0.9U L=0.24U
M14 TP2 AIN GVSS 0 nch W=0.9U L=0.24U
M15 TP1 BIN VDD VDD pch W=1.4U L=0.24U
M16 VDD CIN TP1 VDD pch W=1.4U L=0.24U
M17 TP2 BIN GVSS 0 nch W=0.9U L=0.24U
M18 GVSS CIN TP2 0 nch W=0.9U L=0.24U
M19 VDD AIN TP4 VDD pch W=2.1U L=0.24U
M20 TP4 BIN TP5 VDD pch W=2.1U L=0.24U
M21 TP5 CIN TP3 VDD pch W=2.1U L=0.24U
M22 TP6 CIN TP3 0 nch W=1.3U L=0.24U
M23 TP7 BIN TP6 0 nch W=1.3U L=0.24U
M24 GVSS AIN TP7 0 nch W=1.3U L=0.24U
M26 OUTS TP3 GVSS 0 nch W=0.9U L=0.24U
M28 OUTC TP0 GVSS 0 nch W=1U L=0.24U
M25 OUTS TP3 VDD VDD pch W=1.3U L=0.24U
M27 OUTC TP0 VDD VDD pch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_fadd1s2 OUTS OUTC AIN BIN CIN
M1 TP9 AIN VDD VDD pch W=1.8U L=0.24U
M2 TP0 BIN TP9 VDD pch W=1.7U L=0.24U
M3 TP0 BIN TP8 0 nch W=1.1U L=0.24U
M4 TP8 AIN GVSS 0 nch W=1.2U L=0.24U
M5 TP10 AIN VDD VDD pch W=1.8U L=0.24U
M6 VDD BIN TP10 VDD pch W=1.8U L=0.24U
M7 TP10 CIN TP0 VDD pch W=1.7U L=0.24U
M8 TP11 CIN TP0 0 nch W=1.1U L=0.24U
M9 GVSS BIN TP11 0 nch W=1.2U L=0.24U
M10 TP11 AIN GVSS 0 nch W=1.2U L=0.24U
M11 TP1 AIN VDD VDD pch W=2.1U L=0.24U
M12 TP3 TP0 TP1 VDD pch W=1.66U L=0.24U
M13 TP3 TP0 TP2 0 nch W=1.16U L=0.24U
M14 TP2 AIN GVSS 0 nch W=1.16U L=0.24U
M15 TP1 BIN VDD VDD pch W=2.1U L=0.24U
M16 VDD CIN TP1 VDD pch W=2.1U L=0.24U
M17 TP2 BIN GVSS 0 nch W=1.16U L=0.24U
M18 GVSS CIN TP2 0 nch W=1.16U L=0.24U
M19 VDD AIN TP4 VDD pch W=3.16U L=0.24U
M20 TP4 BIN TP5 VDD pch W=3.16U L=0.24U
M21 TP5 CIN TP3 VDD pch W=3.16U L=0.24U
M22 TP6 CIN TP3 0 nch W=1.74U L=0.24U
M23 TP7 BIN TP6 0 nch W=1.74U L=0.24U
M24 GVSS AIN TP7 0 nch W=1.74U L=0.24U
M26 OUTS TP3 GVSS 0 nch W=1.44U L=0.24U
M28 OUTC TP0 GVSS 0 nch W=1.62U L=0.24U
M25 OUTS TP3 VDD VDD pch W=2.1U L=0.24U
M27 OUTC TP0 VDD VDD pch W=2.32U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_fadd1s3 OUTS OUTC AIN BIN CIN
M1 TP9 AIN VDD VDD pch W=2.7U L=0.24U
M2 TP0 BIN TP9 VDD pch W=2.6U L=0.24U
M3 TP0 BIN TP8 0 nch W=1.6U L=0.24U
M4 TP8 AIN GVSS 0 nch W=1.7U L=0.24U
M5 TP10 AIN VDD VDD pch W=2.7U L=0.24U
M6 VDD BIN TP10 VDD pch W=2.7U L=0.24U
M7 TP10 CIN TP0 VDD pch W=2.6U L=0.24U
M8 TP11 CIN TP0 0 nch W=1.6U L=0.24U
M9 GVSS BIN TP11 0 nch W=1.7U L=0.24U
M10 TP11 AIN GVSS 0 nch W=1.7U L=0.24U
M11 TP1 AIN VDD VDD pch W=2.9U L=0.24U
M12 TP3 TP0 TP1 VDD pch W=2.8U L=0.24U
M13 TP3 TP0 TP2 0 nch W=1.52U L=0.24U
M14 TP2 AIN GVSS 0 nch W=1.52U L=0.24U
M15 TP1 BIN VDD VDD pch W=2.9U L=0.24U
M16 VDD CIN TP1 VDD pch W=2.9U L=0.24U
M17 TP2 BIN GVSS 0 nch W=1.52U L=0.24U
M18 GVSS CIN TP2 0 nch W=1.52U L=0.24U
M19 VDD AIN TP4 VDD pch W=4.4U L=0.24U
M20 TP4 BIN TP5 VDD pch W=4.4U L=0.24U
M21 TP5 CIN TP3 VDD pch W=4.3U L=0.24U
M22 TP6 CIN TP3 0 nch W=2.26U L=0.24U
M23 TP7 BIN TP6 0 nch W=2.26U L=0.24U
M24 GVSS AIN TP7 0 nch W=2.26U L=0.24U
M26 OUTS TP3 GVSS 0 nch W=3.1U L=0.24U
M28 OUTC TP0 GVSS 0 nch W=3.4U L=0.24U
M25 OUTS TP3 VDD VDD pch W=4.2U L=0.24U
M27 OUTC TP0 VDD VDD pch W=4.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_faddpgs1 AIN BIN CIN OUTG OUTP OUTS
M24 OUTG N1N525 GVSS 0 nch W=0.9U L=0.24U
M23 OUTG N1N525 VDD VDD pch W=1.9U L=0.24U
M19 N1N525 AIN N1N553 0 nch W=0.8U L=0.24U
M17 VDD AIN N1N525 VDD pch W=0.9U L=0.24U
M18 N1N525 BIN VDD VDD pch W=0.9U L=0.24U
M20 N1N553 BIN GVSS 0 nch W=0.8U L=0.24U
M5 N1N515 AIN BIN VDD pch W=1.2U L=0.24U
M6 BIN N1N569 N1N515 0 nch W=0.8U L=0.24U
M1 N1N569 AIN VDD VDD pch W=1.5U L=0.24U
M8 BIN AIN N1N623 0 nch W=0.8U L=0.24U
M3 N1N572 CIN VDD VDD pch W=1.5U L=0.24U
M4 N1N572 CIN GVSS 0 nch W=0.7U L=0.24U
M2 N1N569 AIN GVSS 0 nch W=0.7U L=0.24U
M7 N1N623 N1N569 BIN VDD pch W=1.2U L=0.24U
M13 N1N515 BIN AIN VDD pch W=1.6U L=0.24U
M14 N1N515 BIN N1N569 0 nch W=0.7U L=0.24U
M16 N1N623 BIN AIN 0 nch W=0.7U L=0.24U
M15 N1N623 BIN N1N569 VDD pch W=1.6U L=0.24U
M9 N1N693 N1N515 N1N572 VDD pch W=1.2U L=0.24U
M10 N1N572 N1N623 N1N693 0 nch W=0.7U L=0.24U
M11 N1N693 N1N623 CIN VDD pch W=1.2U L=0.24U
M12 CIN N1N515 N1N693 0 nch W=0.7U L=0.24U
M21 OUTS N1N693 VDD VDD pch W=1.4U L=0.24U
M22 OUTS N1N693 GVSS 0 nch W=0.9U L=0.24U
M25 OUTP N1N623 VDD VDD pch W=1.9U L=0.24U
M26 OUTP N1N623 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_faddpgs2 AIN BIN CIN OUTG OUTP OUTS
M24 OUTG N1N525 GVSS 0 nch W=1.1U L=0.24U
M23 OUTG N1N525 VDD VDD pch W=2.47U L=0.24U
M19 N1N525 AIN N1N553 0 nch W=0.96U L=0.24U
M17 VDD AIN N1N525 VDD pch W=1.16U L=0.24U
M18 N1N525 BIN VDD VDD pch W=1.16U L=0.24U
M20 N1N553 BIN GVSS 0 nch W=0.96U L=0.24U
M5 N1N515 AIN BIN VDD pch W=1.56U L=0.24U
M6 BIN N1N569 N1N515 0 nch W=1U L=0.24U
M1 N1N569 AIN VDD VDD pch W=1.96U L=0.24U
M8 BIN AIN N1N623 0 nch W=1U L=0.24U
M3 N1N572 CIN VDD VDD pch W=1.96U L=0.24U
M4 N1N572 CIN GVSS 0 nch W=0.92U L=0.24U
M2 N1N569 AIN GVSS 0 nch W=0.92U L=0.24U
M7 N1N623 N1N569 BIN VDD pch W=1.5U L=0.24U
M13 N1N515 BIN AIN VDD pch W=1.92U L=0.24U
M14 N1N515 BIN N1N569 0 nch W=0.84U L=0.24U
M16 N1N623 BIN AIN 0 nch W=0.84U L=0.24U
M15 N1N623 BIN N1N569 VDD pch W=1.92U L=0.24U
M9 N1N693 N1N515 N1N572 VDD pch W=1.56U L=0.24U
M10 N1N572 N1N623 N1N693 0 nch W=0.84U L=0.24U
M11 N1N693 N1N623 CIN VDD pch W=1.56U L=0.24U
M12 CIN N1N515 N1N693 0 nch W=0.84U L=0.24U
M21 OUTS N1N693 VDD VDD pch W=1.82U L=0.24U
M22 OUTS N1N693 GVSS 0 nch W=1.26U L=0.24U
M25 OUTP N1N623 VDD VDD pch W=2.47U L=0.24U
M26 OUTP N1N623 GVSS 0 nch W=1.68U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_faddpgs3 AIN BIN CIN OUTG OUTP OUTS
M24 OUTG N1N525 GVSS 0 nch W=1.85U L=0.24U
M23 OUTG N1N525 VDD VDD pch W=3.72U L=0.24U
M19 N1N525 AIN N1N553 0 nch W=1.44U L=0.24U
M17 VDD AIN N1N525 VDD pch W=1.74U L=0.24U
M18 N1N525 BIN VDD VDD pch W=1.74U L=0.24U
M20 N1N553 BIN GVSS 0 nch W=1.44U L=0.24U
M5 N1N515 AIN BIN VDD pch W=2.2U L=0.24U
M6 BIN N1N569 N1N515 0 nch W=1.6U L=0.24U
M1 N1N569 AIN VDD VDD pch W=2.94U L=0.24U
M8 BIN AIN N1N623 0 nch W=1.6U L=0.24U
M3 N1N572 CIN VDD VDD pch W=2.34U L=0.24U
M4 N1N572 CIN GVSS 0 nch W=1.18U L=0.24U
M2 N1N569 AIN GVSS 0 nch W=1.38U L=0.24U
M7 N1N623 N1N569 BIN VDD pch W=2.2U L=0.24U
M13 N1N515 BIN AIN VDD pch W=2.92U L=0.24U
M14 N1N515 BIN N1N569 0 nch W=1.3U L=0.24U
M16 N1N623 BIN AIN 0 nch W=1.3U L=0.24U
M15 N1N623 BIN N1N569 VDD pch W=2.92U L=0.24U
M9 N1N693 N1N515 N1N572 VDD pch W=2.34U L=0.24U
M10 N1N572 N1N623 N1N693 0 nch W=1.26U L=0.24U
M11 N1N693 N1N623 CIN VDD pch W=2.34U L=0.24U
M12 CIN N1N515 N1N693 0 nch W=1.26U L=0.24U
M21 OUTS N1N693 VDD VDD pch W=2.7U L=0.24U
M22 OUTS N1N693 GVSS 0 nch W=2.1U L=0.24U
M25 OUTP N1N623 VDD VDD pch W=3.71U L=0.24U
M26 OUTP N1N623 GVSS 0 nch W=2.72U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_hadd1s1 AIN BIN OUTS OUTC
M10 GVSS BIN N1N458 0 nch W=0.7U L=0.24U
M7 N1N450 BIN N1N452 VDD pch W=1.6U L=0.24U
M1 N1N439 AIN VDD VDD pch W=0.8U L=0.24U
M5 N1N452 N1N439 VDD VDD pch W=0.8U L=0.24U
M2 VDD BIN N1N439 VDD pch W=0.8U L=0.24U
M6 VDD AIN N1N450 VDD pch W=1.6U L=0.24U
M3 N1N439 AIN N1N443 0 nch W=0.76U L=0.24U
M4 N1N443 BIN GVSS 0 nch W=0.76U L=0.24U
M8 N1N452 N1N439 N1N458 0 nch W=0.7U L=0.24U
M9 N1N458 AIN GVSS 0 nch W=0.7U L=0.24U
M12 OUTS N1N452 GVSS 0 nch W=1.16U L=0.24U
M14 OUTC N1N439 GVSS 0 nch W=1.4U L=0.24U
M13 OUTC N1N439 VDD VDD pch W=2U L=0.24U
M11 OUTS N1N452 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_hadd1s2 AIN BIN OUTS OUTC
M10 GVSS BIN N1N458 0 nch W=1.1U L=0.24U
M7 N1N450 BIN N1N452 VDD pch W=2.68U L=0.24U
M1 N1N439 AIN VDD VDD pch W=1.4U L=0.24U
M5 N1N452 N1N439 VDD VDD pch W=1.34U L=0.24U
M2 VDD BIN N1N439 VDD pch W=1.4U L=0.24U
M6 VDD AIN N1N450 VDD pch W=2.68U L=0.24U
M3 N1N439 AIN N1N443 0 nch W=1.14U L=0.24U
M4 N1N443 BIN GVSS 0 nch W=1.14U L=0.24U
M8 N1N452 N1N439 N1N458 0 nch W=1.1U L=0.24U
M9 N1N458 AIN GVSS 0 nch W=1.1U L=0.24U
M12 OUTS N1N452 GVSS 0 nch W=1.74U L=0.24U
M14 OUTC N1N439 GVSS 0 nch W=2.1U L=0.24U
M13 OUTC N1N439 VDD VDD pch W=3U L=0.24U
M11 OUTS N1N452 VDD VDD pch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_hadd1s3 AIN BIN OUTS OUTC
M10 GVSS BIN N1N458 0 nch W=2.2U L=0.24U
M7 N1N450 BIN N1N452 VDD pch W=5.6U L=0.24U
M1 N1N439 AIN VDD VDD pch W=2.9U L=0.24U
M5 N1N452 N1N439 VDD VDD pch W=2.8U L=0.24U
M2 VDD BIN N1N439 VDD pch W=2.9U L=0.24U
M6 VDD AIN N1N450 VDD pch W=5.6U L=0.24U
M3 N1N439 AIN N1N443 0 nch W=2.28U L=0.24U
M4 N1N443 BIN GVSS 0 nch W=2.28U L=0.24U
M8 N1N452 N1N439 N1N458 0 nch W=2.2U L=0.24U
M9 N1N458 AIN GVSS 0 nch W=2.2U L=0.24U
M12 OUTS N1N452 GVSS 0 nch W=3.48U L=0.24U
M14 OUTC N1N439 GVSS 0 nch W=4.4U L=0.24U
M13 OUTC N1N439 VDD VDD pch W=6U L=0.24U
M11 OUTS N1N452 VDD VDD pch W=5.94U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_hi1s1 Q DIN
M2 Q DIN GVSS 0 nch W=0.6U L=0.8U
M1 Q DIN VDD VDD pch W=1U L=0.3U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_hib1s1 Q DIN
M2 Q GVSS TP0 VDD pch W=4U L=0.24U
M3 Q VDD TP1 0 nch W=2U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.9U L=0.4U
M4 TP1 DIN GVSS 0 nch W=0.76U L=0.7U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_hnb1s1 Q DIN
M5 Q VDD TP2 0 nch W=2U L=0.24U
M4 Q GVSS TP1 VDD pch W=4U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.6U L=0.24U
M2 TP0 DIN GVSS 0 nch W=0.7U L=0.24U
M3 TP1 TP0 VDD VDD pch W=1.9U L=0.4U
M6 TP2 TP0 GVSS 0 nch W=0.76U L=0.7U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s1 Q DIN
M1 Q DIN VDD VDD pch W=2U L=0.24U
M2 Q DIN GVSS 0 nch W=0.82U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s10 DIN Q
M1 N1N255 DIN VDD VDD pch W=10.5U L=0.24U
M2 N1N255 DIN GVSS 0 nch W=6.8U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=21.8U L=0.24U
M4 N1N266 N1N255 GVSS 0 nch W=13.6U L=0.24U
M5 Q N1N266 VDD VDD pch W=51.6U L=0.24U
M6 Q N1N266 GVSS 0 nch W=20.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s11 DIN Q
M3 N1N255 N1N253 VDD VDD pch W=9U L=0.24U
M4 N1N255 N1N253 GVSS 0 nch W=4.5U L=0.24U
M5 N1N266 N1N255 VDD VDD pch W=20U L=0.24U
M6 N1N266 N1N255 GVSS 0 nch W=11U L=0.24U
M7 N1N268 N1N266 VDD VDD pch W=40U L=0.24U
M8 N1N268 N1N266 GVSS 0 nch W=26U L=0.24U
M1 N1N253 DIN VDD VDD pch W=4U L=0.24U
M2 N1N253 DIN GVSS 0 nch W=2.2U L=0.24U
M9 Q N1N268 VDD VDD pch W=84U L=0.24U
M10 Q N1N268 GVSS 0 nch W=42U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s12 DIN Q
M3 N1N255 N1N253 VDD VDD pch W=16.5U L=0.24U
M4 N1N255 N1N253 GVSS 0 nch W=9.8U L=0.24U
M5 N1N266 N1N255 VDD VDD pch W=36.4U L=0.24U
M6 N1N266 N1N255 GVSS 0 nch W=20.6U L=0.24U
M7 N1N268 N1N266 VDD VDD pch W=88.3U L=0.24U
M8 N1N268 N1N266 GVSS 0 nch W=50.9U L=0.24U
M1 N1N253 DIN VDD VDD pch W=8.3U L=0.24U
M2 N1N253 DIN GVSS 0 nch W=5U L=0.24U
M9 Q N1N268 VDD VDD pch W=180.8U L=0.24U
M10 Q N1N268 GVSS 0 nch W=78.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s2 Q DIN
M1 Q DIN VDD VDD pch W=3.5U L=0.24U
M2 Q DIN GVSS 0 nch W=1.38U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s3 Q DIN
M1 Q DIN VDD VDD pch W=6.22U L=0.24U
M2 Q DIN GVSS 0 nch W=2.68U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s4 Q DIN
M1 Q DIN VDD VDD pch W=7.8U L=0.24U
M2 Q DIN GVSS 0 nch W=3.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s5 Q DIN
M1 Q DIN VDD VDD pch W=9.54U L=0.24U
M2 Q DIN GVSS 0 nch W=4.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s6 Q DIN
M1 Q DIN VDD VDD pch W=12.6U L=0.24U
M2 Q DIN GVSS 0 nch W=5.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s7 Q DIN
M1 N1N255 DIN VDD VDD pch W=4.5U L=0.24U
M2 N1N255 DIN GVSS 0 nch W=2.1U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=5.3U L=0.24U
M4 N1N266 N1N255 GVSS 0 nch W=4U L=0.24U
M5 Q N1N266 VDD VDD pch W=16.5U L=0.24U
M6 Q N1N266 GVSS 0 nch W=9.52U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s8 DIN Q
M1 N1N255 DIN VDD VDD pch W=6.2U L=0.24U
M2 N1N255 DIN GVSS 0 nch W=4.5U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=13.5U L=0.24U
M4 N1N266 N1N255 GVSS 0 nch W=9.5U L=0.24U
M5 Q N1N266 VDD VDD pch W=28.5U L=0.24U
M6 Q N1N266 GVSS 0 nch W=14.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_i1s9 Q DIN
M1 N1N255 DIN VDD VDD pch W=7.3U L=0.24U
M2 N1N255 DIN GVSS 0 nch W=5.2U L=0.24U
M3 N1N266 N1N255 VDD VDD pch W=15.6U L=0.24U
M4 N1N266 N1N255 GVSS 0 nch W=11.2U L=0.24U
M5 Q N1N266 VDD VDD pch W=35.8U L=0.24U
M6 Q N1N266 GVSS 0 nch W=15U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s1 Q DIN
M2 Q DIN GVSS 0 nch W=1.2U L=0.24U
M1 Q DIN VDD VDD pch W=2.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s10 DIN Q
M2 Q DIN GVSS 0 nch W=11.1U L=0.24U
M1 Q DIN VDD VDD pch W=25U L=0.24U
M13 Q DIN VDD VDD pch W=25U L=0.24U
M14 Q DIN GVSS 0 nch W=11.1U L=0.24U
M3 Q DIN VDD VDD pch W=25U L=0.24U
M5 Q DIN VDD VDD pch W=25U L=0.24U
M7 Q DIN VDD VDD pch W=25U L=0.24U
M9 Q DIN VDD VDD pch W=25U L=0.24U
M11 Q DIN VDD VDD pch W=25U L=0.24U
M4 Q DIN GVSS 0 nch W=11.1U L=0.24U
M6 Q DIN GVSS 0 nch W=11.1U L=0.24U
M8 Q DIN GVSS 0 nch W=11.1U L=0.24U
M10 Q DIN GVSS 0 nch W=11.1U L=0.24U
M12 Q DIN GVSS 0 nch W=11.1U L=0.24U
M15 Q DIN VDD VDD pch W=25U L=0.24U
M17 Q DIN VDD VDD pch W=25U L=0.24U
M19 Q DIN VDD VDD pch W=25U L=0.24U
M16 Q DIN GVSS 0 nch W=11.1U L=0.24U
M18 Q DIN GVSS 0 nch W=11.1U L=0.24U
M20 Q DIN GVSS 0 nch W=11.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s11 DIN Q
M2 Q DIN GVSS 0 nch W=23U L=0.24U
M1 Q DIN VDD VDD pch W=50U L=0.24U
M13 Q DIN VDD VDD pch W=50U L=0.24U
M14 Q DIN GVSS 0 nch W=23U L=0.24U
M3 Q DIN VDD VDD pch W=50U L=0.24U
M5 Q DIN VDD VDD pch W=50U L=0.24U
M7 Q DIN VDD VDD pch W=50U L=0.24U
M9 Q DIN VDD VDD pch W=50U L=0.24U
M11 Q DIN VDD VDD pch W=50U L=0.24U
M4 Q DIN GVSS 0 nch W=23U L=0.24U
M6 Q DIN GVSS 0 nch W=23U L=0.24U
M8 Q DIN GVSS 0 nch W=23U L=0.24U
M10 Q DIN GVSS 0 nch W=23U L=0.24U
M12 Q DIN GVSS 0 nch W=23U L=0.24U
M15 Q DIN VDD VDD pch W=50U L=0.24U
M17 Q DIN VDD VDD pch W=50U L=0.24U
M19 Q DIN VDD VDD pch W=50U L=0.24U
M16 Q DIN GVSS 0 nch W=23U L=0.24U
M18 Q DIN GVSS 0 nch W=23U L=0.24U
M20 Q DIN GVSS 0 nch W=23U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s12 DIN Q
M2 Q DIN GVSS 0 nch W=47U L=0.24U
M1 Q DIN VDD VDD pch W=101U L=0.24U
M13 Q DIN VDD VDD pch W=101U L=0.24U
M14 Q DIN GVSS 0 nch W=47U L=0.24U
M3 Q DIN VDD VDD pch W=101U L=0.24U
M5 Q DIN VDD VDD pch W=101U L=0.24U
M7 Q DIN VDD VDD pch W=101U L=0.24U
M9 Q DIN VDD VDD pch W=101U L=0.24U
M11 Q DIN VDD VDD pch W=101U L=0.24U
M4 Q DIN GVSS 0 nch W=47U L=0.24U
M6 Q DIN GVSS 0 nch W=47U L=0.24U
M8 Q DIN GVSS 0 nch W=47U L=0.24U
M10 Q DIN GVSS 0 nch W=47U L=0.24U
M12 Q DIN GVSS 0 nch W=47U L=0.24U
M15 Q DIN VDD VDD pch W=101U L=0.24U
M17 Q DIN VDD VDD pch W=101U L=0.24U
M19 Q DIN VDD VDD pch W=101U L=0.24U
M16 Q DIN GVSS 0 nch W=47U L=0.24U
M18 Q DIN GVSS 0 nch W=47U L=0.24U
M20 Q DIN GVSS 0 nch W=47U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s2 Q DIN
M2 Q DIN GVSS 0 nch W=1.2U L=0.24U
M1 Q DIN VDD VDD pch W=2.9U L=0.24U
M4 Q DIN GVSS 0 nch W=1.2U L=0.24U
M3 Q DIN VDD VDD pch W=2.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s3 Q DIN
M2 Q DIN GVSS 0 nch W=1.2U L=0.24U
M1 Q DIN VDD VDD pch W=2.9U L=0.24U
M4 Q DIN GVSS 0 nch W=1.2U L=0.24U
M3 Q DIN VDD VDD pch W=2.9U L=0.24U
M6 Q DIN GVSS 0 nch W=1.2U L=0.24U
M5 Q DIN VDD VDD pch W=2.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s4 Q DIN
M2 Q DIN GVSS 0 nch W=1.1U L=0.24U
M1 Q DIN VDD VDD pch W=2.6U L=0.24U
M4 Q DIN GVSS 0 nch W=1.1U L=0.24U
M3 Q DIN VDD VDD pch W=2.6U L=0.24U
M6 Q DIN GVSS 0 nch W=1.1U L=0.24U
M5 Q DIN VDD VDD pch W=2.6U L=0.24U
M7 Q DIN VDD VDD pch W=2.6U L=0.24U
M8 Q DIN GVSS 0 nch W=1.1U L=0.24U
M10 Q DIN GVSS 0 nch W=1.1U L=0.24U
M9 Q DIN VDD VDD pch W=2.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s5 Q DIN
M2 Q DIN GVSS 0 nch W=1.1U L=0.24U
M1 Q DIN VDD VDD pch W=2.5U L=0.24U
M4 Q DIN GVSS 0 nch W=1.1U L=0.24U
M3 Q DIN VDD VDD pch W=2.5U L=0.24U
M6 Q DIN GVSS 0 nch W=1.1U L=0.24U
M5 Q DIN VDD VDD pch W=2.5U L=0.24U
M7 Q DIN VDD VDD pch W=2.5U L=0.24U
M8 Q DIN GVSS 0 nch W=1.1U L=0.24U
M10 Q DIN GVSS 0 nch W=1.1U L=0.24U
M9 Q DIN VDD VDD pch W=2.5U L=0.24U
M12 Q DIN GVSS 0 nch W=1.1U L=0.24U
M11 Q DIN VDD VDD pch W=2.5U L=0.24U
M14 Q DIN GVSS 0 nch W=1.1U L=0.24U
M13 Q DIN VDD VDD pch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s6 DIN Q
M2 Q DIN GVSS 0 nch W=1.1U L=0.24U
M1 Q DIN VDD VDD pch W=2.5U L=0.24U
M4 Q DIN GVSS 0 nch W=1.1U L=0.24U
M3 Q DIN VDD VDD pch W=2.5U L=0.24U
M6 Q DIN GVSS 0 nch W=1.1U L=0.24U
M5 Q DIN VDD VDD pch W=2.5U L=0.24U
M7 Q DIN VDD VDD pch W=2.5U L=0.24U
M8 Q DIN GVSS 0 nch W=1.1U L=0.24U
M10 Q DIN GVSS 0 nch W=1.1U L=0.24U
M9 Q DIN VDD VDD pch W=2.5U L=0.24U
M12 Q DIN GVSS 0 nch W=1.1U L=0.24U
M11 Q DIN VDD VDD pch W=2.5U L=0.24U
M19 Q DIN VDD VDD pch W=2.5U L=0.24U
M13 Q DIN VDD VDD pch W=2.5U L=0.24U
M16 Q DIN GVSS 0 nch W=1.1U L=0.24U
M18 Q DIN GVSS 0 nch W=1.1U L=0.24U
M17 Q DIN VDD VDD pch W=2.5U L=0.24U
M14 Q DIN GVSS 0 nch W=1.1U L=0.24U
M15 Q DIN VDD VDD pch W=2.5U L=0.24U
M20 Q DIN GVSS 0 nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s7 DIN Q
M2 Q DIN GVSS 0 nch W=1.8U L=0.24U
M1 Q DIN VDD VDD pch W=4.2U L=0.24U
M13 Q DIN VDD VDD pch W=4.2U L=0.24U
M14 Q DIN GVSS 0 nch W=1.8U L=0.24U
M3 Q DIN VDD VDD pch W=4.2U L=0.24U
M5 Q DIN VDD VDD pch W=4.2U L=0.24U
M7 Q DIN VDD VDD pch W=4.2U L=0.24U
M9 Q DIN VDD VDD pch W=4.2U L=0.24U
M11 Q DIN VDD VDD pch W=4.2U L=0.24U
M4 Q DIN GVSS 0 nch W=1.8U L=0.24U
M6 Q DIN GVSS 0 nch W=1.8U L=0.24U
M8 Q DIN GVSS 0 nch W=1.8U L=0.24U
M10 Q DIN GVSS 0 nch W=1.8U L=0.24U
M12 Q DIN GVSS 0 nch W=1.8U L=0.24U
M15 Q DIN VDD VDD pch W=4.2U L=0.24U
M17 Q DIN VDD VDD pch W=4.2U L=0.24U
M19 Q DIN VDD VDD pch W=4.2U L=0.24U
M16 Q DIN GVSS 0 nch W=1.8U L=0.24U
M18 Q DIN GVSS 0 nch W=1.8U L=0.24U
M20 Q DIN GVSS 0 nch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s8 DIN Q
M2 Q DIN GVSS 0 nch W=3.2U L=0.24U
M1 Q DIN VDD VDD pch W=7.5U L=0.24U
M13 Q DIN VDD VDD pch W=7.5U L=0.24U
M14 Q DIN GVSS 0 nch W=3.2U L=0.24U
M3 Q DIN VDD VDD pch W=7.5U L=0.24U
M5 Q DIN VDD VDD pch W=7.5U L=0.24U
M7 Q DIN VDD VDD pch W=7.5U L=0.24U
M9 Q DIN VDD VDD pch W=7.5U L=0.24U
M11 Q DIN VDD VDD pch W=7.5U L=0.24U
M4 Q DIN GVSS 0 nch W=3.2U L=0.24U
M6 Q DIN GVSS 0 nch W=3.2U L=0.24U
M8 Q DIN GVSS 0 nch W=3.2U L=0.24U
M10 Q DIN GVSS 0 nch W=3.2U L=0.24U
M12 Q DIN GVSS 0 nch W=3.2U L=0.24U
M15 Q DIN VDD VDD pch W=7.5U L=0.24U
M17 Q DIN VDD VDD pch W=7.5U L=0.24U
M19 Q DIN VDD VDD pch W=7.5U L=0.24U
M16 Q DIN GVSS 0 nch W=3.2U L=0.24U
M18 Q DIN GVSS 0 nch W=3.2U L=0.24U
M20 Q DIN GVSS 0 nch W=3.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ib1s9 DIN Q
M2 Q DIN GVSS 0 nch W=6U L=0.24U
M1 Q DIN VDD VDD pch W=14U L=0.24U
M13 Q DIN VDD VDD pch W=14U L=0.24U
M14 Q DIN GVSS 0 nch W=6U L=0.24U
M3 Q DIN VDD VDD pch W=14U L=0.24U
M5 Q DIN VDD VDD pch W=14U L=0.24U
M7 Q DIN VDD VDD pch W=14U L=0.24U
M9 Q DIN VDD VDD pch W=14U L=0.24U
M11 Q DIN VDD VDD pch W=14U L=0.24U
M4 Q DIN GVSS 0 nch W=6U L=0.24U
M6 Q DIN GVSS 0 nch W=6U L=0.24U
M8 Q DIN GVSS 0 nch W=6U L=0.24U
M10 Q DIN GVSS 0 nch W=6U L=0.24U
M12 Q DIN GVSS 0 nch W=6U L=0.24U
M15 Q DIN VDD VDD pch W=14U L=0.24U
M17 Q DIN VDD VDD pch W=14U L=0.24U
M19 Q DIN VDD VDD pch W=14U L=0.24U
M16 Q DIN GVSS 0 nch W=6U L=0.24U
M18 Q DIN GVSS 0 nch W=6U L=0.24U
M20 Q DIN GVSS 0 nch W=6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lclks1 DIN CLK QN Q
M10 QN TP1 GVSS 0 nch W=1.56U L=0.24U
M4 TP1 TP0 DIN VDD pch W=1.8U L=0.24U
M3 DIN CLK TP1 0 nch W=0.8U L=0.24U
M8 TP2 QN GVSS 0 nch W=0.8U L=0.24U
M11 Q QN VDD VDD pch W=2.92U L=0.24U
M12 Q QN GVSS 0 nch W=1.34U L=0.24U
M9 QN TP1 VDD VDD pch W=2.92U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M6 TP1 TP0 TP2 0 nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lclks2 DIN CLK QN Q
M10 QN TP1 GVSS 0 nch W=3.38U L=0.24U
M4 TP1 TP0 DIN VDD pch W=2.2U L=0.24U
M3 DIN CLK TP1 0 nch W=1U L=0.24U
M8 TP2 QN GVSS 0 nch W=0.8U L=0.24U
M11 Q QN VDD VDD pch W=6.06U L=0.24U
M12 Q QN GVSS 0 nch W=2.88U L=0.24U
M9 QN TP1 VDD VDD pch W=6.16U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M6 TP1 TP0 TP2 0 nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lcs1 CLRB DIN CLK QN Q
M9 QN TP1 VDD VDD pch W=3.1U L=0.24U
M10 QN CLRB VDD VDD pch W=3.1U L=0.24U
M12 TP3 CLRB GVSS 0 nch W=2.56U L=0.24U
M11 QN TP1 TP3 0 nch W=2.56U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK GVSS 0 nch W=0.8U L=0.24U
M4 TP1 TP0 DIN VDD pch W=1.88U L=0.24U
M3 DIN CLK TP1 0 nch W=0.84U L=0.24U
M6 TP1 TP0 TP2 0 nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M8 TP2 QN GVSS 0 nch W=0.8U L=0.24U
M13 Q QN VDD VDD pch W=3.16U L=0.24U
M14 Q QN GVSS 0 nch W=1.48U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lcs2 CLRB DIN CLK QN Q
M9 QN TP1 VDD VDD pch W=5.6U L=0.24U
M10 QN CLRB VDD VDD pch W=5.6U L=0.24U
M12 TP3 CLRB GVSS 0 nch W=5.1U L=0.24U
M11 QN TP1 TP3 0 nch W=5.1U L=0.24U
M1 TP0 CLK VDD VDD pch W=1.3U L=0.24U
M2 TP0 CLK GVSS 0 nch W=0.8U L=0.24U
M4 TP1 TP0 DIN VDD pch W=2.38U L=0.24U
M3 DIN CLK TP1 0 nch W=1.56U L=0.24U
M6 TP1 TP0 TP2 0 nch W=0.8U L=0.24U
M5 TP2 CLK TP1 VDD pch W=1.8U L=0.24U
M7 TP2 QN VDD VDD pch W=1.3U L=0.24U
M8 TP2 QN GVSS 0 nch W=0.8U L=0.24U
M13 Q QN VDD VDD pch W=6.36U L=0.24U
M14 Q QN GVSS 0 nch W=2.94U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lnnds1 Q QN SIN RIN
M1 Q SIN  VDD  VDD P  W=1.56u   L=0.24U
M2 Q QN VDD  VDD P  W=1.56u   L=0.24U
M3 Q QN TP0  GVSS   N  W=1.02U   L=0.24U
M4 TP0 SIN  GVSS    GVSS   N  W=1.02u   L=0.24U
M5 VDD Q  QN VDD P  W=1.56u   L=0.24U
M6 VDD RIN  QN VDD P  W=1.56u   L=0.24U
M7 TP1 Q  QN GVSS   N  W=1.02U   L=0.24U
M8 GVSS   RIN  TP1  GVSS   N  W=1.02u   L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lnnds2 Q QN SIN RIN
M1 Q SIN  VDD  VDD P  W=3.16u  L=0.24U
M2 Q QN VDD  VDD P  W=3.16u  L=0.24U
M3 Q QN TP0  GVSS   N  W=2.06U  L=0.24U
M4 TP0 SIN  GVSS    GVSS   N  W=2.06u  L=0.24U
M5 VDD Q  QN VDD P  W=3.16u  L=0.24U
M6 VDD RIN  QN VDD P  W=3.16u  L=0.24U
M7 TP1 Q  QN GVSS   N  W=2.06U  L=0.24U
M8 GVSS   RIN  TP1  GVSS   N  W=2.06u  L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lnors1 Q QN RIN SIN
M1  TP0   SIN   VDD    VDD  pch W=3.54u    L=0.24U
M2  QN  Q   TP0    VDD  pch W=3.54u    L=0.24U
M3  QN  SIN   GVSS      GVSS    nch W=0.9u     L=0.24U
M4  GVSS     Q   QN   GVSS    nch W=0.9u     L=0.24U
M5  VDD  RIN    TP1    VDD  pch W=3.54u    L=0.24U
M6  TP1  QN   Q    VDD  pch W=3.54u    L=0.24U
M7  Q  QN   GVSS      GVSS    nch W=0.9u     L=0.24U
M8  GVSS    RIN    Q    GVSS    nch W=0.9u     L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lnors2 Q QN RIN SIN
M1  TP0   SIN   VDD    VDD  pch W=7.18u    L=0.24U
M2  QN  Q   TP0    VDD  pch W=7.18u    L=0.24U
M3  QN  SIN   GVSS      GVSS    nch W=1.8u     L=0.24U
M4  GVSS     Q   QN   GVSS    nch W=1.8u     L=0.24U
M5  VDD  RIN    TP1    VDD  pch W=7.18u    L=0.24U
M6  TP1  QN   Q    VDD  pch W=7.18u    L=0.24U
M7  Q  QN   GVSS      GVSS    nch W=1.8u     L=0.24U
M8  GVSS    RIN    Q    GVSS    nch W=1.8u     L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lscs1 CLK DIN SETB CLRB QN Q
M18 Q TP5 GVSS 0 nch W=1.88U L=0.24U
M11 TP5 TP4 TP2 VDD pch W=1.8U L=0.24U
M12 TP2 CLK TP5 0 nch W=1.3U L=0.24U
M16 TP6 Q GVSS 0 nch W=0.8U L=0.24U
M19 QN Q VDD VDD pch W=2.96U L=0.24U
M20 QN Q GVSS 0 nch W=1.32U L=0.24U
M17 Q TP5 VDD VDD pch W=2.98U L=0.24U
M15 TP6 Q VDD VDD pch W=1.3U L=0.24U
M13 TP5 TP4 TP6 0 nch W=0.8U L=0.24U
M14 TP6 CLK TP5 VDD pch W=1.8U L=0.24U
M9 TP4 CLK VDD VDD pch W=1.3U L=0.24U
M10 TP4 CLK GVSS 0 nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
M5 TP2 CLRB VDD VDD pch W=2U L=0.24U
M4 TP2 DIN TP1 VDD pch W=2U L=0.24U
M6 TP2 CLRB TP3 0 nch W=1U L=0.24U
M7 TP3 DIN GVSS 0 nch W=1U L=0.24U
M8 TP3 TP0 GVSS 0 nch W=1U L=0.24U
M3 TP1 TP0 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lscs2 CLK DIN SETB CLRB QN Q
M18 Q TP5 GVSS 0 nch W=3.98U L=0.24U
M11 TP5 TP4 TP2 VDD pch W=2.8U L=0.24U
M12 TP2 CLK TP5 0 nch W=2.6U L=0.24U
M16 TP6 Q GVSS 0 nch W=0.8U L=0.24U
M19 QN Q VDD VDD pch W=5.96U L=0.24U
M20 QN Q GVSS 0 nch W=2.42U L=0.24U
M17 Q TP5 VDD VDD pch W=6.02U L=0.24U
M15 TP6 Q VDD VDD pch W=1.3U L=0.24U
M13 TP5 TP4 TP6 0 nch W=0.8U L=0.24U
M14 TP6 CLK TP5 VDD pch W=1.3U L=0.24U
M9 TP4 CLK VDD VDD pch W=1.3U L=0.24U
M10 TP4 CLK GVSS 0 nch W=0.8U L=0.24U
M1 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M2 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
M5 TP2 CLRB VDD VDD pch W=2.5U L=0.24U
M4 TP2 DIN TP1 VDD pch W=2.5U L=0.24U
M6 TP2 CLRB TP3 0 nch W=1.3U L=0.24U
M7 TP3 DIN GVSS 0 nch W=1.3U L=0.24U
M8 TP3 TP0 GVSS 0 nch W=1.3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lss1 SETB DIN CLK QN Q
M11 Q TP2 VDD VDD pch W=3.14U L=0.24U
M12 Q SETB VDD VDD pch W=3.14U L=0.24U
M14 TP4 SETB GVSS 0 nch W=2.88U L=0.24U
M13 Q TP2 TP4 0 nch W=2.88U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M4 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M6 TP2 TP1 TP0 VDD pch W=2.2U L=0.24U
M5 TP0 CLK TP2 0 nch W=1.8U L=0.24U
M8 TP2 TP1 TP3 0 nch W=0.8U L=0.24U
M7 TP3 CLK TP2 VDD pch W=1.3U L=0.24U
M9 TP3 Q VDD VDD pch W=1.3U L=0.24U
M10 TP3 Q GVSS 0 nch W=0.8U L=0.24U
M15 QN Q VDD VDD pch W=3.12U L=0.24U
M16 QN Q GVSS 0 nch W=1.4U L=0.24U
M2 TP0 DIN GVSS 0 nch W=0.9U L=0.24U
M1 TP0 DIN VDD VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_lss2 SETB DIN CLK QN Q
M11 Q TP2 VDD VDD pch W=6.9U L=0.24U
M12 Q SETB VDD VDD pch W=6.9U L=0.24U
M14 TP4 SETB GVSS 0 nch W=6.6U L=0.24U
M13 Q TP2 TP4 0 nch W=6.6U L=0.24U
M3 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M4 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M6 TP2 TP1 TP0 VDD pch W=2.8U L=0.24U
M5 TP0 CLK TP2 0 nch W=2.5U L=0.24U
M8 TP2 TP1 TP3 0 nch W=0.8U L=0.24U
M7 TP3 CLK TP2 VDD pch W=1.3U L=0.24U
M9 TP3 Q VDD VDD pch W=1.3U L=0.24U
M10 TP3 Q GVSS 0 nch W=0.8U L=0.24U
M15 QN Q VDD VDD pch W=6.8U L=0.24U
M16 QN Q GVSS 0 nch W=3U L=0.24U
M2 TP0 DIN GVSS 0 nch W=1.42U L=0.24U
M1 TP0 DIN VDD VDD pch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mx21s1 Q DIN1 SIN DIN2
M4 DIN2 SIN N1N438 0 nch W=0.6U L=0.24U
M3 N1N438 N1N434 DIN1 0 nch W=0.6U L=0.24U
M2 N1N434 SIN GVSS 0 nch W=0.6U L=0.24U
M1 N1N434 SIN VDD VDD pch W=1.2U L=0.24U
M7 N1N441 N1N438 GVSS 0 nch W=1U L=0.24U
M9 Q N1N441 GVSS 0 nch W=1U L=0.24U
M6 N1N441 N1N438 VDD VDD pch W=1.3U L=0.24U
M8 Q N1N441 VDD VDD pch W=2.4U L=0.24U
M5 N1N438 N1N441 VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mx21s2 Q DIN1 SIN DIN2
M4 DIN2 SIN N1N438 0 nch W=0.6U L=0.24U
M3 N1N438 N1N430 DIN2 VDD pch W=1.1U L=0.24U
M7 N1N498 N1N438 VDD VDD pch W=1.6U L=0.24U
M8 N1N498 N1N438 GVSS 0 nch W=0.7U L=0.24U
M2 DIN1 N1N430 N1N438 0 nch W=0.6U L=0.24U
M1 N1N438 SIN DIN1 VDD pch W=1.1U L=0.24U
M6 N1N430 SIN GVSS 0 nch W=0.7U L=0.24U
M5 N1N430 SIN VDD VDD pch W=1.4U L=0.24U
M9 Q N1N498 VDD VDD pch W=3U L=0.24U
M10 Q N1N498 GVSS 0 nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mx21s3 Q DIN1 SIN DIN2
M6 N1N430 SIN GVSS 0 nch W=0.9U L=0.24U
M5 N1N430 SIN VDD VDD pch W=1.8U L=0.24U
M3 N1N438 N1N430 DIN2 VDD pch W=1.8U L=0.24U
M4 DIN2 SIN N1N438 0 nch W=0.9U L=0.24U
M2 DIN1 N1N430 N1N438 0 nch W=0.9U L=0.24U
M1 N1N438 SIN DIN1 VDD pch W=1.8U L=0.24U
M8 N1N483 N1N438 GVSS 0 nch W=0.9U L=0.24U
M10 Q N1N483 GVSS 0 nch W=3.6U L=0.24U
M7 N1N483 N1N438 VDD VDD pch W=2.2U L=0.24U
M9 Q N1N483 VDD VDD pch W=5.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mx41s1 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M3 N1N440 N1N429 DIN1 0 nch W=0.8U L=0.24U
M4 N1N440 SIN0 DIN2 0 nch W=0.8U L=0.24U
M5 N1N442 N1N429 DIN3 0 nch W=0.8U L=0.24U
M6 N1N442 SIN0 DIN4 0 nch W=0.8U L=0.24U
M10 N1N448 SIN1 N1N442 0 nch W=0.6U L=0.24U
M9 N1N448 N1N451 N1N440 0 nch W=0.6U L=0.24U
M2 N1N429 SIN0 GVSS 0 nch W=0.6U L=0.24U
M1 N1N429 SIN0 VDD VDD pch W=1.2U L=0.24U
M7 N1N451 SIN1 VDD VDD pch W=1.2U L=0.24U
M8 N1N451 SIN1 GVSS 0 nch W=0.6U L=0.24U
M13 N1N458 N1N448 GVSS 0 nch W=1.1U L=0.24U
M12 N1N458 N1N448 VDD VDD pch W=2U L=0.24U
M14 Q N1N458 VDD VDD pch W=2.5U L=0.24U
M15 Q N1N458 GVSS 0 nch W=1.3U L=0.24U
M11 N1N448 N1N458 VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mx41s2 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M2 DIN1 N1N564 N1N488 0 nch W=0.8U L=0.24U
M1 N1N488 SIN0 DIN1 VDD pch W=1.6U L=0.24U
M3 N1N488 N1N564 DIN2 VDD pch W=1.6U L=0.24U
M4 DIN2 SIN0 N1N488 0 nch W=0.8U L=0.24U
M5 N1N490 SIN0 DIN3 VDD pch W=1.6U L=0.24U
M6 DIN3 N1N564 N1N490 0 nch W=0.8U L=0.24U
M7 N1N490 N1N564 DIN4 VDD pch W=1.6U L=0.24U
M8 DIN4 SIN0 N1N490 0 nch W=0.8U L=0.24U
M10 N1N564 SIN0 GVSS 0 nch W=0.8U L=0.24U
M9 N1N564 SIN0 VDD VDD pch W=1.6U L=0.24U
M11 N1N507 SIN1 VDD VDD pch W=1.2U L=0.24U
M12 N1N507 SIN1 GVSS 0 nch W=0.6U L=0.24U
M15 N1N510 N1N507 N1N490 VDD pch W=1.2U L=0.24U
M16 N1N490 SIN1 N1N510 0 nch W=0.6U L=0.24U
M13 N1N510 SIN1 N1N488 VDD pch W=1.2U L=0.24U
M14 N1N488 N1N507 N1N510 0 nch W=0.6U L=0.24U
M17 N1N646 N1N510 VDD VDD pch W=2.4U L=0.24U
M19 Q N1N646 VDD VDD pch W=3.3U L=0.24U
M18 N1N646 N1N510 GVSS 0 nch W=1U L=0.24U
M20 Q N1N646 GVSS 0 nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mx41s3 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M14 N1N490 SIN1 N1N510 0 nch W=0.9U L=0.24U
M13 N1N510 N1N507 N1N490 VDD pch W=1.8U L=0.24U
M2 DIN1 N1N493 N1N488 0 nch W=1.2U L=0.24U
M1 N1N488 SIN0 DIN1 VDD pch W=2.4U L=0.24U
M4 DIN2 SIN0 N1N488 0 nch W=1.2U L=0.24U
M3 N1N488 N1N493 DIN2 VDD pch W=2.4U L=0.24U
M5 N1N490 SIN0 DIN3 VDD pch W=2.4U L=0.24U
M6 DIN3 N1N493 N1N490 0 nch W=1.2U L=0.24U
M7 N1N490 N1N493 DIN4 VDD pch W=2.4U L=0.24U
M8 DIN4 SIN0 N1N490 0 nch W=1.2U L=0.24U
M11 N1N510 SIN1 N1N488 VDD pch W=1.8U L=0.24U
M12 N1N488 N1N507 N1N510 0 nch W=0.9U L=0.24U
M17 Q N1N569 VDD VDD pch W=6.6U L=0.24U
M18 Q N1N569 GVSS 0 nch W=4U L=0.24U
M10 N1N493 SIN0 GVSS 0 nch W=1.2U L=0.24U
M9 N1N493 SIN0 VDD VDD pch W=2.5U L=0.24U
M19 N1N507 SIN1 VDD VDD pch W=1.8U L=0.24U
M20 N1N507 SIN1 GVSS 0 nch W=0.9U L=0.24U
M15 N1N569 N1N510 VDD VDD pch W=3.5U L=0.24U
M16 N1N569 N1N510 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mxi21s1 Q DIN1 SIN DIN2
M4 DIN2 SIN N1N438 0 nch W=0.6U L=0.24U
M7 Q N1N438 GVSS 0 nch W=2.4U L=0.24U
M6 Q N1N438 VDD VDD pch W=2.4U L=0.24U
M1 N1N434 SIN VDD VDD pch W=1.2U L=0.24U
M2 N1N434 SIN GVSS 0 nch W=0.6U L=0.24U
M3 N1N438 N1N434 DIN1 0 nch W=0.6U L=0.24U
M5 N1N438 Q VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mxi21s2 Q DIN1 SIN DIN2
M8 Q N1N438 GVSS 0 nch W=1.24U L=0.24U
M6 DIN2 SIN N1N438 0 nch W=0.6U L=0.24U
M7 Q N1N438 VDD VDD pch W=3U L=0.24U
M5 N1N438 N1N430 DIN2 VDD pch W=1.1U L=0.24U
M4 DIN1 N1N430 N1N438 0 nch W=0.6U L=0.24U
M3 N1N438 SIN DIN1 VDD pch W=1.1U L=0.24U
M2 N1N430 SIN GVSS 0 nch W=0.7U L=0.24U
M1 N1N430 SIN VDD VDD pch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mxi21s3 Q DIN1 SIN DIN2
M8 Q N1N438 GVSS 0 nch W=2.1U L=0.24U
M6 DIN2 SIN N1N438 0 nch W=0.9U L=0.24U
M7 Q N1N438 VDD VDD pch W=5.7U L=0.24U
M5 N1N438 N1N430 DIN2 VDD pch W=1.8U L=0.24U
M4 DIN1 N1N430 N1N438 0 nch W=0.9U L=0.24U
M3 N1N438 SIN DIN1 VDD pch W=1.8U L=0.24U
M2 N1N430 SIN GVSS 0 nch W=0.9U L=0.24U
M1 N1N430 SIN VDD VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mxi41s1 Q DIN1 SIN0 SIN1 DIN2 DIN3 DIN4
M3 N1N440 N1N429 DIN1 0 nch W=0.8U L=0.24U
M4 N1N440 SIN0 DIN2 0 nch W=0.8U L=0.24U
M5 N1N442 N1N429 DIN3 0 nch W=0.8U L=0.24U
M6 N1N442 SIN0 DIN4 0 nch W=0.8U L=0.24U
M10 N1N448 SIN1 N1N442 0 nch W=0.6U L=0.24U
M9 N1N448 N1N451 N1N440 0 nch W=0.6U L=0.24U
M13 Q N1N448 GVSS 0 nch W=1.7U L=0.24U
M12 Q N1N448 VDD VDD pch W=2.5U L=0.24U
M2 N1N429 SIN0 GVSS 0 nch W=0.6U L=0.24U
M1 N1N429 SIN0 VDD VDD pch W=1.2U L=0.24U
M8 N1N451 SIN1 GVSS 0 nch W=0.6U L=0.24U
M7 N1N451 SIN1 VDD VDD pch W=1.2U L=0.24U
M11 N1N448 Q VDD VDD pch W=0.6U L=0.4U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mxi41s2 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M18 Q N1N510 GVSS 0 nch W=1.5U L=0.24U
M16 N1N490 SIN1 N1N510 0 nch W=0.6U L=0.24U
M15 N1N510 N1N589 N1N490 VDD pch W=1.2U L=0.24U
M17 Q N1N510 VDD VDD pch W=3.4U L=0.24U
M2 DIN1 N1N493 N1N488 0 nch W=0.8U L=0.24U
M1 N1N488 SIN0 DIN1 VDD pch W=1.6U L=0.24U
M4 DIN2 SIN0 N1N488 0 nch W=0.8U L=0.24U
M3 N1N488 N1N493 DIN2 VDD pch W=1.6U L=0.24U
M6 DIN3 N1N493 N1N490 0 nch W=0.8U L=0.24U
M5 N1N490 SIN0 DIN3 VDD pch W=1.6U L=0.24U
M8 DIN4 SIN0 N1N490 0 nch W=0.8U L=0.24U
M7 N1N490 N1N493 DIN4 VDD pch W=1.6U L=0.24U
M9 N1N493 SIN0 VDD VDD pch W=1.6U L=0.24U
M10 N1N493 SIN0 GVSS 0 nch W=0.8U L=0.24U
M11 N1N589 SIN1 VDD VDD pch W=1.2U L=0.24U
M12 N1N589 SIN1 GVSS 0 nch W=0.6U L=0.24U
M14 N1N488 N1N589 N1N510 0 nch W=0.6U L=0.24U
M13 N1N510 SIN1 N1N488 VDD pch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_mxi41s3 Q DIN1 SIN1 SIN0 DIN2 DIN3 DIN4
M18 Q N1N510 GVSS 0 nch W=2.2U L=0.24U
M16 N1N490 SIN1 N1N510 0 nch W=0.9U L=0.24U
M15 N1N510 N1N589 N1N490 VDD pch W=1.8U L=0.24U
M17 Q N1N510 VDD VDD pch W=5.7U L=0.24U
M2 DIN1 N1N493 N1N488 0 nch W=1.2U L=0.24U
M1 N1N488 SIN0 DIN1 VDD pch W=2.4U L=0.24U
M4 DIN2 SIN0 N1N488 0 nch W=1.2U L=0.24U
M3 N1N488 N1N493 DIN2 VDD pch W=2.4U L=0.24U
M6 DIN3 N1N493 N1N490 0 nch W=1.2U L=0.24U
M5 N1N490 SIN0 DIN3 VDD pch W=2.4U L=0.24U
M8 DIN4 SIN0 N1N490 0 nch W=1.2U L=0.24U
M7 N1N490 N1N493 DIN4 VDD pch W=2.4U L=0.24U
M9 N1N493 SIN0 VDD VDD pch W=2.5U L=0.24U
M10 N1N493 SIN0 GVSS 0 nch W=1.2U L=0.24U
M11 N1N589 SIN1 VDD VDD pch W=1.8U L=0.24U
M12 N1N589 SIN1 GVSS 0 nch W=0.9U L=0.24U
M14 N1N488 N1N589 N1N510 0 nch W=0.9U L=0.24U
M13 N1N510 SIN1 N1N488 VDD pch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s1 Q DIN
M4 Q N1N262 GVSS 0 nch W=1.5U L=0.24U
M3 Q N1N262 VDD VDD pch W=2.5U L=0.24U
M1 N1N262 DIN VDD VDD pch W=2.1U L=0.24U
M2 N1N262 DIN GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s10 Q DIN
M4 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M3 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M1 N1N318 DIN VDD VDD pch W=43U L=0.24U
M2 N1N318 DIN GVSS 0 nch W=20U L=0.24U
M6 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M5 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M7 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M8 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M10 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M9 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M11 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M12 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M14 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M13 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M15 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M16 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s11 DIN Q
M4 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M3 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M1 N1N318 DIN VDD VDD pch W=53U L=0.24U
M2 N1N318 DIN GVSS 0 nch W=24U L=0.24U
M6 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M5 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M7 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M8 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M10 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M9 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M11 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M12 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M14 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
M13 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M15 Q N1N318 VDD VDD pch W=6.6U L=0.24U
M16 Q N1N318 GVSS 0 nch W=3.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s12 DIN Q
M4 Q N1N318 GVSS 0 nch W=3.7U L=0.24U
M3 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M1 N1N318 DIN VDD VDD pch W=55U L=0.24U
M2 N1N318 DIN GVSS 0 nch W=27U L=0.24U
M6 Q N1N318 GVSS 0 nch W=3.7U L=0.24U
M5 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M7 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M8 Q N1N318 GVSS 0 nch W=3.7U L=0.24U
M10 Q N1N318 GVSS 0 nch W=3.7U L=0.24U
M9 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M11 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M12 Q N1N318 GVSS 0 nch W=3.7U L=0.24U
M14 Q N1N318 GVSS 0 nch W=3.7U L=0.24U
M13 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M15 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M16 Q N1N318 GVSS 0 nch W=3.7U L=0.24U
M17 Q N1N318 VDD VDD pch W=6.5U L=0.24U
M18 Q N1N318 GVSS 0 nch W=3.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s2 Q DIN
M4 Q N1N262 GVSS 0 nch W=1.5U L=0.24U
M3 Q N1N262 VDD VDD pch W=2.8U L=0.24U
M1 N1N262 DIN VDD VDD pch W=2.5U L=0.24U
M2 N1N262 DIN GVSS 0 nch W=1.4U L=0.24U
M6 Q N1N262 GVSS 0 nch W=1.5U L=0.24U
M5 Q N1N262 VDD VDD pch W=2.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s3 Q DIN
M4 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M3 Q N1N262 VDD VDD pch W=2.3U L=0.24U
M1 N1N262 DIN VDD VDD pch W=3.9U L=0.24U
M2 N1N262 DIN GVSS 0 nch W=1.6U L=0.24U
M6 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M5 Q N1N262 VDD VDD pch W=2.3U L=0.24U
M7 Q N1N262 VDD VDD pch W=2.3U L=0.24U
M8 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s4 Q DIN
M4 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M3 Q N1N262 VDD VDD pch W=2U L=0.24U
M1 N1N262 DIN VDD VDD pch W=4U L=0.24U
M2 N1N262 DIN GVSS 0 nch W=2U L=0.24U
M6 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M5 Q N1N262 VDD VDD pch W=2U L=0.24U
M7 Q N1N262 VDD VDD pch W=2U L=0.24U
M8 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M10 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M9 Q N1N262 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s5 Q DIN
M4 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M3 Q N1N262 VDD VDD pch W=2U L=0.24U
M1 N1N262 DIN VDD VDD pch W=5.5U L=0.24U
M2 N1N262 DIN GVSS 0 nch W=2.6U L=0.24U
M6 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M5 Q N1N262 VDD VDD pch W=2U L=0.24U
M7 Q N1N262 VDD VDD pch W=2U L=0.24U
M8 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M10 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
M9 Q N1N262 VDD VDD pch W=2U L=0.24U
M11 Q N1N262 VDD VDD pch W=2U L=0.24U
M12 Q N1N262 GVSS 0 nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s6 Q DIN
M4 Q N1N318 GVSS 0 nch W=1.1U L=0.24U
M3 Q N1N318 VDD VDD pch W=2U L=0.24U
M1 N1N318 DIN VDD VDD pch W=6.2U L=0.24U
M2 N1N318 DIN GVSS 0 nch W=3U L=0.24U
M6 Q N1N318 GVSS 0 nch W=1.1U L=0.24U
M5 Q N1N318 VDD VDD pch W=2U L=0.24U
M7 Q N1N318 VDD VDD pch W=2U L=0.24U
M8 Q N1N318 GVSS 0 nch W=1.1U L=0.24U
M10 Q N1N318 GVSS 0 nch W=1.1U L=0.24U
M9 Q N1N318 VDD VDD pch W=2U L=0.24U
M11 Q N1N318 VDD VDD pch W=2U L=0.24U
M12 Q N1N318 GVSS 0 nch W=1.1U L=0.24U
M14 Q N1N318 GVSS 0 nch W=1.1U L=0.24U
M13 Q N1N318 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s7 DIN Q
M4 Q N1N318 GVSS 0 nch W=1.7U L=0.24U
M3 Q N1N318 VDD VDD pch W=3U L=0.24U
M1 N1N318 DIN VDD VDD pch W=8U L=0.24U
M2 N1N318 DIN GVSS 0 nch W=3.8U L=0.24U
M6 Q N1N318 GVSS 0 nch W=1.7U L=0.24U
M5 Q N1N318 VDD VDD pch W=3U L=0.24U
M7 Q N1N318 VDD VDD pch W=3U L=0.24U
M8 Q N1N318 GVSS 0 nch W=1.7U L=0.24U
M10 Q N1N318 GVSS 0 nch W=1.7U L=0.24U
M9 Q N1N318 VDD VDD pch W=3U L=0.24U
M11 Q N1N318 VDD VDD pch W=3U L=0.24U
M12 Q N1N318 GVSS 0 nch W=1.7U L=0.24U
M14 Q N1N318 GVSS 0 nch W=1.7U L=0.24U
M13 Q N1N318 VDD VDD pch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s8 DIN Q
M4 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M3 Q N1N318 VDD VDD pch W=4U L=0.24U
M1 N1N318 DIN VDD VDD pch W=15U L=0.24U
M2 N1N318 DIN GVSS 0 nch W=7U L=0.24U
M6 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M5 Q N1N318 VDD VDD pch W=4U L=0.24U
M7 Q N1N318 VDD VDD pch W=4U L=0.24U
M8 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M10 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M9 Q N1N318 VDD VDD pch W=4U L=0.24U
M11 Q N1N318 VDD VDD pch W=4U L=0.24U
M12 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M14 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M13 Q N1N318 VDD VDD pch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nb1s9 DIN Q
M4 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M3 Q N1N318 VDD VDD pch W=4U L=0.24U
M1 N1N318 DIN VDD VDD pch W=26U L=0.24U
M2 N1N318 DIN GVSS 0 nch W=12U L=0.24U
M6 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M5 Q N1N318 VDD VDD pch W=4U L=0.24U
M7 Q N1N318 VDD VDD pch W=4U L=0.24U
M8 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M10 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M9 Q N1N318 VDD VDD pch W=4U L=0.24U
M11 Q N1N318 VDD VDD pch W=4U L=0.24U
M12 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M14 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
M13 Q N1N318 VDD VDD pch W=4U L=0.24U
M15 Q N1N318 VDD VDD pch W=4U L=0.24U
M16 Q N1N318 GVSS 0 nch W=2.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd2s1 Q DIN1 DIN2
M3 Q DIN1 N1N275 0 nch W=1.16U L=0.24U
M1 Q DIN1 VDD VDD pch W=1.8U L=0.24U
M2 VDD DIN2 Q VDD pch W=1.8U L=0.24U
M4 N1N275 DIN2 GVSS 0 nch W=1.16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd2s2 Q DIN1 DIN2
M3 Q DIN1 N1N275 0 nch W=2.18U L=0.24U
M1 Q DIN1 VDD VDD pch W=3.3U L=0.24U
M2 VDD DIN2 Q VDD pch W=3.3U L=0.24U
M4 N1N275 DIN2 GVSS 0 nch W=2.18U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd2s3 Q DIN1 DIN2
M3 Q DIN1 N1N275 0 nch W=4U L=0.24U
M1 Q DIN1 VDD VDD pch W=5.9U L=0.24U
M2 VDD DIN2 Q VDD pch W=5.9U L=0.24U
M4 N1N275 DIN2 GVSS 0 nch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd3s1 Q DIN1 DIN2 DIN3
M4 Q DIN1 N1N260 0 nch W=1.5U L=0.24U
M3 Q DIN3 VDD VDD pch W=1.8U L=0.24U
M2 Q DIN2 VDD VDD pch W=1.8U L=0.24U
M1 Q DIN1 VDD VDD pch W=1.8U L=0.24U
M6 N1N293 DIN3 GVSS 0 nch W=1.5U L=0.24U
M5 N1N260 DIN2 N1N293 0 nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd3s2 Q DIN1 DIN2 DIN3
M4 Q DIN1 N1N260 0 nch W=2.64U L=0.24U
M3 Q DIN3 VDD VDD pch W=3.12U L=0.24U
M2 Q DIN2 VDD VDD pch W=3.12U L=0.24U
M1 Q DIN1 VDD VDD pch W=3.12U L=0.24U
M6 N1N293 DIN3 GVSS 0 nch W=2.64U L=0.24U
M5 N1N260 DIN2 N1N293 0 nch W=2.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd3s3 Q DIN1 DIN2 DIN3
M4 Q DIN1 N1N260 0 nch W=4.8U L=0.24U
M3 Q DIN3 VDD VDD pch W=6U L=0.24U
M2 Q DIN2 VDD VDD pch W=6U L=0.24U
M1 Q DIN1 VDD VDD pch W=6U L=0.24U
M6 N1N293 DIN3 GVSS 0 nch W=5.6U L=0.24U
M5 N1N260 DIN2 N1N293 0 nch W=5.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd4s1 Q DIN1 DIN2 DIN3 DIN4
M1 Q DIN1 VDD VDD pch W=1.9U L=0.24U
M2 Q DIN2 VDD VDD pch W=1.9U L=0.24U
M3 Q DIN3 VDD VDD pch W=1.9U L=0.24U
M4 Q DIN4 VDD VDD pch W=1.9U L=0.24U
M5 Q DIN1 N1N348 0 nch W=1.8U L=0.24U
M6 N1N348 DIN2 N1N347 0 nch W=1.84U L=0.24U
M7 N1N347 DIN3 N1N346 0 nch W=1.94U L=0.24U
M8 N1N346 DIN4 GVSS 0 nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd4s2 Q DIN1 DIN2 DIN3 DIN4
M1 Q DIN1 VDD VDD pch W=3.12U L=0.24U
M2 Q DIN2 VDD VDD pch W=3.12U L=0.24U
M3 Q DIN3 VDD VDD pch W=3.12U L=0.24U
M4 Q DIN4 VDD VDD pch W=3.12U L=0.24U
M5 Q DIN1 N1N348 0 nch W=2.98U L=0.24U
M6 N1N348 DIN2 N1N347 0 nch W=3U L=0.24U
M7 N1N347 DIN3 N1N346 0 nch W=3.1U L=0.24U
M8 N1N346 DIN4 GVSS 0 nch W=3.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd4s3 Q DIN1 DIN2 DIN3 DIN4
M4 N1N280 DIN2 GVSS 0 nch W=4.1U L=0.24U
M3 N1N269 DIN1 N1N280 0 nch W=3.1U L=0.24U
M14 Q N1N315 GVSS 0 nch W=4U L=0.24U
M12 GVSS N1N298 N1N315 0 nch W=3.1U L=0.24U
M11 N1N315 N1N269 GVSS 0 nch W=3.1U L=0.24U
M8 N1N309 DIN4 GVSS 0 nch W=4.1U L=0.24U
M7 N1N298 DIN3 N1N309 0 nch W=3.1U L=0.24U
M5 N1N298 DIN3 VDD VDD pch W=3.7U L=0.24U
M6 VDD DIN4 N1N298 VDD pch W=3.7U L=0.24U
M10 N1N325 N1N298 N1N315 VDD pch W=7.2U L=0.24U
M1 N1N269 DIN1 VDD VDD pch W=3.7U L=0.24U
M2 VDD DIN2 N1N269 VDD pch W=3.7U L=0.24U
M9 N1N325 N1N269 VDD VDD pch W=7.5U L=0.24U
M13 Q N1N315 VDD VDD pch W=8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd5s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M4 N1N442 DIN1 N1N438 0 nch W=3.9U L=0.24U
M1 N1N442 DIN1 VDD VDD pch W=4.2U L=0.24U
M2 N1N442 DIN2 VDD VDD pch W=4.2U L=0.24U
M3 N1N442 DIN3 VDD VDD pch W=4.2U L=0.24U
M5 N1N438 DIN2 N1N440 0 nch W=4.8U L=0.24U
M6 N1N440 DIN3 GVSS 0 nch W=5.8U L=0.24U
M11 N1N446 N1N442 VDD VDD pch W=6.7U L=0.24U
M12 N1N446 N1N455 N1N448 VDD pch W=6.1U L=0.24U
M13 N1N448 N1N442 GVSS 0 nch W=3.1U L=0.24U
M14 GVSS N1N455 N1N448 0 nch W=3.1U L=0.24U
M7 N1N455 DIN4 VDD VDD pch W=4.2U L=0.24U
M8 N1N455 DIN5 VDD VDD pch W=4.2U L=0.24U
M9 N1N455 DIN4 N1N457 0 nch W=3.4U L=0.24U
M10 N1N457 DIN5 GVSS 0 nch W=3.9U L=0.24U
M15 Q N1N448 VDD VDD pch W=4.3U L=0.24U
M16 Q N1N448 GVSS 0 nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd6s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M1 N1N419 DIN1 VDD VDD pch W=4.1U L=0.24U
M2 N1N419 DIN2 VDD VDD pch W=4.1U L=0.24U
M3 N1N419 DIN3 VDD VDD pch W=4.1U L=0.24U
M4 N1N419 DIN1 N1N429 0 nch W=3.9U L=0.24U
M5 N1N429 DIN2 N1N428 0 nch W=4.8U L=0.24U
M6 N1N428 DIN3 GVSS 0 nch W=5.8U L=0.24U
M13 N1N427 N1N419 VDD VDD pch W=6.7U L=0.24U
M14 N1N427 N1N424 N1N425 VDD pch W=6.1U L=0.24U
M15 N1N425 N1N419 GVSS 0 nch W=3U L=0.24U
M16 GVSS N1N424 N1N425 0 nch W=3U L=0.24U
M10 N1N424 DIN4 N1N453 0 nch W=3.9U L=0.24U
M7 N1N424 DIN4 VDD VDD pch W=4.1U L=0.24U
M8 N1N424 DIN5 VDD VDD pch W=4.1U L=0.24U
M9 N1N424 DIN6 VDD VDD pch W=4.1U L=0.24U
M11 N1N453 DIN5 N1N455 0 nch W=4.8U L=0.24U
M12 N1N455 DIN6 GVSS 0 nch W=5.8U L=0.24U
M18 Q N1N425 GVSS 0 nch W=2.1U L=0.24U
M17 Q N1N425 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd7s3 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M1 N1N439 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N439 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 VDD DIN3 N1N439 VDD pch W=2.1U L=0.24U
M4 N1N439 DIN1 N1N425 0 nch W=2.4U L=0.24U
M5 N1N425 DIN2 N1N424 0 nch W=2.6U L=0.24U
M6 N1N424 DIN3 GVSS 0 nch W=2.8U L=0.24U
M11 N1N448 DIN7 VDD VDD pch W=2.1U L=0.24U
M12 N1N448 DIN6 VDD VDD pch W=2.1U L=0.24U
M13 VDD DIN5 N1N448 VDD pch W=2.1U L=0.24U
M14 VDD DIN4 N1N448 VDD pch W=2.1U L=0.24U
M15 N1N448 DIN4 N1N423 0 nch W=6.3U L=0.24U
M16 N1N423 DIN5 N1N422 0 nch W=6.5U L=0.24U
M17 N1N422 DIN6 N1N421 0 nch W=6.7U L=0.24U
M18 N1N421 DIN7 GVSS 0 nch W=6.9U L=0.24U
M7 N1N454 N1N439 VDD VDD pch W=5.2U L=0.24U
M8 N1N454 N1N448 N1N455 VDD pch W=5.2U L=0.24U
M9 N1N455 N1N439 GVSS 0 nch W=2.3U L=0.24U
M10 GVSS N1N448 N1N455 0 nch W=2.3U L=0.24U
M20 Q N1N455 GVSS 0 nch W=2.4U L=0.24U
M19 Q N1N455 VDD VDD pch W=6.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nnd8s3 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 Q
M5 N1N304 DIN1 N1N314 0 nch W=6.3U L=0.24U
M1 N1N304 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N304 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 N1N304 DIN3 VDD VDD pch W=2.1U L=0.24U
M4 N1N304 DIN4 VDD VDD pch W=2.1U L=0.24U
M6 N1N314 DIN2 N1N316 0 nch W=6.5U L=0.24U
M7 N1N316 DIN3 N1N318 0 nch W=6.7U L=0.24U
M8 N1N318 DIN4 GVSS 0 nch W=6.9U L=0.24U
M9 N1N343 N1N304 VDD VDD pch W=5.4U L=0.24U
M10 N1N343 N1N413 N1N345 VDD pch W=5.4U L=0.24U
M11 N1N345 N1N304 GVSS 0 nch W=1.5U L=0.24U
M12 GVSS N1N413 N1N345 0 nch W=1.5U L=0.24U
M13 N1N413 DIN5 VDD VDD pch W=2.1U L=0.24U
M14 N1N413 DIN6 VDD VDD pch W=2.1U L=0.24U
M15 N1N413 DIN7 VDD VDD pch W=2.1U L=0.24U
M16 N1N413 DIN8 VDD VDD pch W=2.1U L=0.24U
M17 N1N413 DIN5 N1N362 0 nch W=6.3U L=0.24U
M18 N1N362 DIN6 N1N364 0 nch W=6.5U L=0.24U
M19 N1N364 DIN7 N1N366 0 nch W=6.7U L=0.24U
M20 N1N366 DIN8 GVSS 0 nch W=6.9U L=0.24U
M22 Q N1N345 GVSS 0 nch W=3U L=0.24U
M21 Q N1N345 VDD VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor2s1 Q DIN1 DIN2
M3 Q DIN1 GVSS 0 nch W=0.7U L=0.24U
M1 N1N427 DIN1 VDD VDD pch W=3U L=0.24U
M2 Q DIN2 N1N427 VDD pch W=3U L=0.24U
M4 Q DIN2 GVSS 0 nch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor2s2 Q DIN1 DIN2
M3 Q DIN1 GVSS 0 nch W=1.5U L=0.24U
M1 N1N427 DIN1 VDD VDD pch W=6.34U L=0.24U
M2 Q DIN2 N1N427 VDD pch W=6.34U L=0.24U
M4 Q DIN2 GVSS 0 nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor2s3 Q DIN1 DIN2
M3 Q DIN1 GVSS 0 nch W=2.7U L=0.24U
M1 N1N427 DIN1 VDD VDD pch W=10.9U L=0.24U
M2 Q DIN2 N1N427 VDD pch W=10.9U L=0.24U
M4 Q DIN2 GVSS 0 nch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor3s1 Q DIN1 DIN2 DIN3
M4 Q DIN1 GVSS 0 nch W=0.74U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=4.38U L=0.24U
M2 N1N430 DIN2 N1N428 VDD pch W=4.38U L=0.24U
M3 Q DIN3 N1N430 VDD pch W=4.38U L=0.24U
M5 Q DIN2 GVSS 0 nch W=0.74U L=0.24U
M6 Q DIN3 GVSS 0 nch W=0.74U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor3s2 Q DIN1 DIN2 DIN3
M4 Q DIN1 GVSS 0 nch W=1.7U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=9.4U L=0.24U
M2 N1N430 DIN2 N1N428 VDD pch W=9.4U L=0.24U
M3 Q DIN3 N1N430 VDD pch W=9.4U L=0.24U
M5 Q DIN2 GVSS 0 nch W=1.7U L=0.24U
M6 Q DIN3 GVSS 0 nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor3s3 Q DIN1 DIN2 DIN3
M4 Q DIN1 GVSS 0 nch W=3.1U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=16U L=0.24U
M2 N1N430 DIN2 N1N428 VDD pch W=16U L=0.24U
M3 Q DIN3 N1N430 VDD pch W=16U L=0.24U
M5 Q DIN2 GVSS 0 nch W=3.1U L=0.24U
M6 Q DIN3 GVSS 0 nch W=3.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor4s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 GVSS 0 nch W=0.86U L=0.24U
M1 N1N452 DIN1 VDD VDD pch W=6.2U L=0.24U
M2 N1N450 DIN2 N1N452 VDD pch W=6U L=0.24U
M3 N1N448 DIN3 N1N450 VDD pch W=5.8U L=0.24U
M4 Q DIN4 N1N448 VDD pch W=5.5U L=0.24U
M6 Q DIN2 GVSS 0 nch W=0.86U L=0.24U
M7 Q DIN3 GVSS 0 nch W=0.86U L=0.24U
M8 Q DIN4 GVSS 0 nch W=0.86U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor4s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 GVSS 0 nch W=1.7U L=0.24U
M1 N1N452 DIN1 VDD VDD pch W=12U L=0.24U
M2 N1N450 DIN2 N1N452 VDD pch W=11.8U L=0.24U
M3 N1N448 DIN3 N1N450 VDD pch W=11.4U L=0.24U
M4 Q DIN4 N1N448 VDD pch W=10.6U L=0.24U
M6 Q DIN2 GVSS 0 nch W=1.7U L=0.24U
M7 Q DIN3 GVSS 0 nch W=1.7U L=0.24U
M8 Q DIN4 GVSS 0 nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor4s3 Q DIN1 DIN2 DIN3 DIN4
M3 N1N438 DIN1 GVSS 0 nch W=1.8U L=0.24U
M1 N1N436 DIN1 VDD VDD pch W=5.2U L=0.24U
M2 N1N438 DIN2 N1N436 VDD pch W=4.4U L=0.24U
M4 N1N438 DIN2 GVSS 0 nch W=1.8U L=0.24U
M5 N1N450 N1N438 VDD VDD pch W=4.2U L=0.24U
M6 VDD N1N457 N1N450 VDD pch W=3.8U L=0.24U
M7 N1N450 N1N438 N1N453 0 nch W=4.4U L=0.24U
M8 N1N453 N1N457 GVSS 0 nch W=4.4U L=0.24U
M9 N1N455 DIN3 VDD VDD pch W=5.2U L=0.24U
M10 N1N457 DIN4 N1N455 VDD pch W=4.4U L=0.24U
M11 N1N457 DIN3 GVSS 0 nch W=1.8U L=0.24U
M12 N1N457 DIN4 GVSS 0 nch W=1.8U L=0.24U
M14 Q N1N450 GVSS 0 nch W=4.2U L=0.24U
M13 Q N1N450 VDD VDD pch W=8.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor5s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 GVSS 0 nch W=0.7U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=3.1U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=2.8U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=2.5U L=0.24U
M4 N1N444 DIN3 GVSS 0 nch W=0.7U L=0.24U
M6 N1N444 DIN1 GVSS 0 nch W=0.7U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=1.9U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=1.7U L=0.24U
M9 N1N494 DIN5 GVSS 0 nch W=0.7U L=0.24U
M10 GVSS DIN4 N1N494 0 nch W=0.7U L=0.24U
M11 N1N474 N1N444 VDD VDD pch W=2U L=0.24U
M12 VDD N1N494 N1N474 VDD pch W=2U L=0.24U
M13 N1N474 N1N444 N1N480 0 nch W=1.6U L=0.24U
M14 N1N480 N1N494 GVSS 0 nch W=1.6U L=0.24U
M16 Q N1N474 GVSS 0 nch W=1.1U L=0.24U
M15 Q N1N474 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor5s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 GVSS 0 nch W=1.4U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=6.1U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=5.9U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=5.7U L=0.24U
M4 N1N444 DIN3 GVSS 0 nch W=1.4U L=0.24U
M6 N1N444 DIN1 GVSS 0 nch W=1.4U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=4U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=3.8U L=0.24U
M9 N1N494 DIN5 GVSS 0 nch W=1.4U L=0.24U
M10 GVSS DIN4 N1N494 0 nch W=1.4U L=0.24U
M11 N1N474 N1N444 VDD VDD pch W=3.9U L=0.24U
M12 VDD N1N494 N1N474 VDD pch W=3.9U L=0.24U
M13 N1N474 N1N444 N1N480 0 nch W=3.7U L=0.24U
M14 N1N480 N1N494 GVSS 0 nch W=3.8U L=0.24U
M16 Q N1N474 GVSS 0 nch W=2.1U L=0.24U
M15 Q N1N474 VDD VDD pch W=4.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor5s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 GVSS 0 nch W=2.3U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=10.7U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=10.2U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=9.5U L=0.24U
M4 N1N444 DIN3 GVSS 0 nch W=2.3U L=0.24U
M6 N1N444 DIN1 GVSS 0 nch W=2.3U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=6.3U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=6.2U L=0.24U
M9 N1N494 DIN5 GVSS 0 nch W=2.3U L=0.24U
M10 GVSS DIN4 N1N494 0 nch W=2.3U L=0.24U
M11 N1N474 N1N444 VDD VDD pch W=6.8U L=0.24U
M12 VDD N1N494 N1N474 VDD pch W=6.8U L=0.24U
M13 N1N474 N1N444 N1N480 0 nch W=5.8U L=0.24U
M14 N1N480 N1N494 GVSS 0 nch W=5.9U L=0.24U
M16 Q N1N474 GVSS 0 nch W=4U L=0.24U
M15 Q N1N474 VDD VDD pch W=8.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor6s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M3 N1N421 DIN3 N1N425 VDD pch W=2.5U L=0.24U
M2 N1N425 DIN2 N1N426 VDD pch W=2.8U L=0.24U
M4 N1N421 DIN3 GVSS 0 nch W=0.7U L=0.24U
M1 N1N426 DIN1 VDD VDD pch W=3.1U L=0.24U
M5 N1N421 DIN2 GVSS 0 nch W=0.7U L=0.24U
M6 N1N421 DIN1 GVSS 0 nch W=0.7U L=0.24U
M11 N1N428 DIN4 VDD VDD pch W=3.1U L=0.24U
M12 N1N423 DIN5 N1N428 VDD pch W=2.8U L=0.24U
M13 N1N434 DIN6 N1N423 VDD pch W=2.5U L=0.24U
M14 N1N434 DIN6 GVSS 0 nch W=0.7U L=0.24U
M8 VDD N1N434 N1N453 VDD pch W=2U L=0.24U
M9 N1N453 N1N421 N1N451 0 nch W=1.6U L=0.24U
M10 N1N451 N1N434 GVSS 0 nch W=1.6U L=0.24U
M16 N1N434 DIN4 GVSS 0 nch W=0.7U L=0.24U
M15 N1N434 DIN5 GVSS 0 nch W=0.7U L=0.24U
M7 N1N453 N1N421 VDD VDD pch W=2U L=0.24U
M18 Q N1N453 GVSS 0 nch W=1.1U L=0.24U
M17 Q N1N453 VDD VDD pch W=2.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor6s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N444 DIN3 GVSS 0 nch W=1.4U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=6.1U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=5.9U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=5.7U L=0.24U
M11 N1N460 DIN4 VDD VDD pch W=6.1U L=0.24U
M5 N1N444 DIN2 GVSS 0 nch W=1.4U L=0.24U
M6 N1N444 DIN1 GVSS 0 nch W=1.4U L=0.24U
M12 N1N462 DIN5 N1N460 VDD pch W=5.9U L=0.24U
M13 N1N464 DIN6 N1N462 VDD pch W=5.7U L=0.24U
M14 N1N464 DIN6 GVSS 0 nch W=1.4U L=0.24U
M15 N1N464 DIN5 GVSS 0 nch W=1.4U L=0.24U
M16 N1N464 DIN4 GVSS 0 nch W=1.4U L=0.24U
M7 N1N480 N1N444 VDD VDD pch W=3.9U L=0.24U
M8 VDD N1N464 N1N480 VDD pch W=3.9U L=0.24U
M9 N1N480 N1N444 N1N483 0 nch W=3.7U L=0.24U
M10 N1N483 N1N464 GVSS 0 nch W=3.8U L=0.24U
M18 Q N1N480 GVSS 0 nch W=2.1U L=0.24U
M17 Q N1N480 VDD VDD pch W=4.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor6s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M4 N1N506 DIN3 GVSS 0 nch W=2.3U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=10.7U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=10.2U L=0.24U
M3 N1N506 DIN3 N1N442 VDD pch W=9.5U L=0.24U
M11 N1N460 DIN4 VDD VDD pch W=10.7U L=0.24U
M5 N1N506 DIN2 GVSS 0 nch W=2.3U L=0.24U
M6 N1N506 DIN1 GVSS 0 nch W=2.3U L=0.24U
M12 N1N462 DIN5 N1N460 VDD pch W=10.2U L=0.24U
M13 N1N464 DIN6 N1N462 VDD pch W=9.5U L=0.24U
M14 N1N464 DIN6 GVSS 0 nch W=2.3U L=0.24U
M15 N1N464 DIN5 GVSS 0 nch W=2.3U L=0.24U
M16 N1N464 DIN4 GVSS 0 nch W=2.3U L=0.24U
M7 N1N480 N1N506 VDD VDD pch W=6.8U L=0.24U
M8 VDD N1N464 N1N480 VDD pch W=6.8U L=0.24U
M9 N1N480 N1N506 N1N483 0 nch W=5.8U L=0.24U
M10 N1N483 N1N464 GVSS 0 nch W=5.9U L=0.24U
M18 Q N1N480 GVSS 0 nch W=4U L=0.24U
M17 Q N1N480 VDD VDD pch W=8.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_nor7s3 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M4 N1N446 DIN1 GVSS 0 nch W=2.34U L=0.24U
M1 N1N441 DIN1 VDD VDD pch W=9U L=0.24U
M2 N1N443 DIN2 N1N441 VDD pch W=8.8U L=0.24U
M3 N1N446 DIN3 N1N443 VDD pch W=8.6U L=0.24U
M5 N1N446 DIN2 GVSS 0 nch W=2.34U L=0.24U
M6 N1N446 DIN3 GVSS 0 nch W=2.34U L=0.24U
M7 N1N465 N1N446 VDD VDD pch W=5.4U L=0.24U
M8 VDD N1N471 N1N465 VDD pch W=5.4U L=0.24U
M9 N1N465 N1N446 N1N473 0 nch W=5U L=0.24U
M10 GVSS N1N471 N1N473 0 nch W=5U L=0.24U
M11 N1N478 DIN4 VDD VDD pch W=11.7U L=0.24U
M12 N1N480 DIN5 N1N478 VDD pch W=11.5U L=0.24U
M13 N1N491 DIN6 N1N480 VDD pch W=11.3U L=0.24U
M16 N1N471 DIN6 GVSS 0 nch W=2.34U L=0.24U
M17 N1N471 DIN5 GVSS 0 nch W=2.34U L=0.24U
M18 N1N471 DIN4 GVSS 0 nch W=2.34U L=0.24U
M15 N1N471 DIN7 GVSS 0 nch W=2.34U L=0.24U
M14 N1N471 DIN7 N1N491 VDD pch W=11.1U L=0.24U
M19 Q N1N465 VDD VDD pch W=7U L=0.24U
M20 Q N1N465 GVSS 0 nch W=3.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_npd1s1 OUTD GIN
M1 OUTD GIN GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_npd1s2 OUTD GIN
M1 OUTD GIN GVSS 0 nch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_npt1s1 DIN OUTD OUTS
M1 OUTD DIN OUTS 0 nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_npt1s2 DIN OUTD OUTS
M1 OUTD DIN OUTS 0 nch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_npt1s3 DIN OUTD OUTS
M1 OUTD DIN OUTS 0 nch W=8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_npt1s4 DIN OUTD OUTS
M1 OUTD DIN OUTS 0 nch W=16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_npt1s5 DIN OUTD OUTS
M1 OUTD DIN OUTS 0 nch W=32U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_npt1s6 DIN OUTS OUTD
M1 OUTD DIN OUTS 0 nch W=65U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oaaoi1123s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 Q DIN7 GVSS 0 nch W=0.6U L=0.24U
M7 Q DIN7 N1N349 VDD pch W=6.9U L=0.24U
M4 N1N349 DIN6 N1N360 VDD pch W=6.9U L=0.24U
M5 N1N360 DIN4 N1N283 VDD pch W=6.9U L=0.24U
M6 N1N349 DIN5 N1N283 VDD pch W=6.9U L=0.24U
M3 VDD DIN3 N1N360 VDD pch W=6.9U L=0.24U
M1 N1N360 DIN2 VDD VDD pch W=6.9U L=0.24U
M2 N1N360 DIN1 VDD VDD pch W=6.9U L=0.24U
M9 Q DIN6 N1N315 0 nch W=1U L=0.24U
M10 N1N289 DIN3 Q 0 nch W=1.3U L=0.24U
M12 N1N315 DIN5 GVSS 0 nch W=1U L=0.24U
M11 N1N315 DIN4 GVSS 0 nch W=1U L=0.24U
M13 N1N289 DIN2 N1N291 0 nch W=1.3U L=0.24U
M14 N1N291 DIN1 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oaaoi1123s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 N1N302 DIN7 GVSS 0 nch W=0.6U L=0.24U
M7 N1N302 DIN7 N1N349 VDD pch W=6.9U L=0.24U
M4 N1N349 DIN6 N1N360 VDD pch W=6.9U L=0.24U
M5 N1N360 DIN4 N1N283 VDD pch W=6.9U L=0.24U
M6 N1N349 DIN5 N1N283 VDD pch W=6.9U L=0.24U
M3 VDD DIN3 N1N360 VDD pch W=6.9U L=0.24U
M1 N1N360 DIN2 VDD VDD pch W=6.9U L=0.24U
M2 N1N360 DIN1 VDD VDD pch W=6.9U L=0.24U
M9 N1N302 DIN6 N1N315 0 nch W=1U L=0.24U
M10 N1N289 DIN3 N1N302 0 nch W=1.3U L=0.24U
M12 N1N315 DIN5 GVSS 0 nch W=1U L=0.24U
M11 N1N315 DIN4 GVSS 0 nch W=1U L=0.24U
M13 N1N289 DIN2 N1N291 0 nch W=1.3U L=0.24U
M14 N1N291 DIN1 GVSS 0 nch W=1.3U L=0.24U
M15 N1N371 N1N302 VDD VDD pch W=3.7U L=0.24U
M16 N1N371 N1N302 GVSS 0 nch W=1.6U L=0.24U
M18 Q N1N371 GVSS 0 nch W=4.1U L=0.24U
M17 Q N1N371 VDD VDD pch W=7.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oaaoi1123s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7
M8 N1N302 DIN7 GVSS 0 nch W=0.6U L=0.24U
M7 N1N302 DIN7 N1N349 VDD pch W=6.9U L=0.24U
M4 N1N349 DIN6 N1N360 VDD pch W=6.9U L=0.24U
M5 N1N360 DIN4 N1N283 VDD pch W=6.9U L=0.24U
M6 N1N349 DIN5 N1N283 VDD pch W=6.9U L=0.24U
M3 VDD DIN3 N1N360 VDD pch W=6.9U L=0.24U
M1 N1N360 DIN2 VDD VDD pch W=6.9U L=0.24U
M2 N1N360 DIN1 VDD VDD pch W=6.9U L=0.24U
M9 N1N302 DIN6 N1N315 0 nch W=1U L=0.24U
M10 N1N289 DIN3 N1N302 0 nch W=1.3U L=0.24U
M12 N1N315 DIN5 GVSS 0 nch W=1U L=0.24U
M11 N1N315 DIN4 GVSS 0 nch W=1U L=0.24U
M13 N1N289 DIN2 N1N291 0 nch W=1.3U L=0.24U
M14 N1N291 DIN1 GVSS 0 nch W=1.3U L=0.24U
M15 N1N371 N1N302 VDD VDD pch W=5.2U L=0.24U
M16 N1N371 N1N302 GVSS 0 nch W=2.2U L=0.24U
M18 Q N1N371 GVSS 0 nch W=5.7U L=0.24U
M17 Q N1N371 VDD VDD pch W=10.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai1112s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N284 0 nch W=1.4U L=0.24U
M1 Q DIN1 VDD VDD pch W=0.7U L=0.24U
M2 Q DIN2 VDD VDD pch W=0.7U L=0.24U
M3 Q DIN3 VDD VDD pch W=0.7U L=0.24U
M4 VDD DIN4 N1N302 VDD pch W=1.4U L=0.24U
M5 N1N302 DIN5 Q VDD pch W=1.4U L=0.24U
M7 N1N284 DIN2 N1N286 0 nch W=1.4U L=0.24U
M8 N1N286 DIN3 N1N292 0 nch W=1.4U L=0.24U
M9 N1N292 DIN4 GVSS 0 nch W=1.4U L=0.24U
M10 GVSS DIN5 N1N292 0 nch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai1112s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN1 N1N284 0 nch W=2U L=0.24U
M1 Q DIN1 VDD VDD pch W=1U L=0.24U
M2 Q DIN2 VDD VDD pch W=1U L=0.24U
M3 Q DIN3 VDD VDD pch W=1U L=0.24U
M4 VDD DIN4 N1N302 VDD pch W=2U L=0.24U
M5 N1N302 DIN5 Q VDD pch W=2U L=0.24U
M7 N1N284 DIN2 N1N286 0 nch W=2U L=0.24U
M8 N1N286 DIN3 N1N292 0 nch W=2U L=0.24U
M9 N1N292 DIN4 GVSS 0 nch W=2U L=0.24U
M10 GVSS DIN5 N1N292 0 nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai1112s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N278 DIN1 N1N284 0 nch W=1.8U L=0.24U
M1 N1N278 DIN1 VDD VDD pch W=0.9U L=0.24U
M2 N1N278 DIN2 VDD VDD pch W=0.9U L=0.24U
M3 N1N278 DIN3 VDD VDD pch W=0.9U L=0.24U
M4 VDD DIN4 N1N302 VDD pch W=1.8U L=0.24U
M5 N1N302 DIN5 N1N278 VDD pch W=1.8U L=0.24U
M7 N1N284 DIN2 N1N286 0 nch W=1.8U L=0.24U
M8 N1N286 DIN3 N1N292 0 nch W=1.9U L=0.24U
M9 N1N292 DIN4 GVSS 0 nch W=1.9U L=0.24U
M10 GVSS DIN5 N1N292 0 nch W=1.9U L=0.24U
M11 N1N326 N1N278 VDD VDD pch W=3.4U L=0.24U
M12 N1N326 N1N278 GVSS 0 nch W=1.8U L=0.24U
M14 Q N1N326 GVSS 0 nch W=3.1U L=0.24U
M13 Q N1N326 VDD VDD pch W=5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai13s1 Q DIN1 DIN2 DIN3 DIN4
M1 N1N330 DIN2 VDD VDD pch W=1.8U L=0.24U
M6 N1N339 DIN2 GVSS 0 nch W=0.7U L=0.24U
M2 N1N332 DIN3 N1N330 VDD pch W=1.8U L=0.24U
M3 Q DIN4 N1N332 VDD pch W=1.8U L=0.24U
M4 VDD DIN1 Q VDD pch W=0.66U L=0.24U
M7 N1N339 DIN3 GVSS 0 nch W=0.7U L=0.24U
M8 GVSS DIN4 N1N339 0 nch W=0.7U L=0.24U
M5 N1N339 DIN1 Q 0 nch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai13s2 Q DIN1 DIN2 DIN3 DIN4
M1 N1N330 DIN2 VDD VDD pch W=2.16U L=0.24U
M6 N1N339 DIN2 GVSS 0 nch W=0.84U L=0.24U
M2 N1N332 DIN3 N1N330 VDD pch W=2.16U L=0.24U
M3 Q DIN4 N1N332 VDD pch W=2.16U L=0.24U
M4 VDD DIN1 Q VDD pch W=0.8U L=0.24U
M7 N1N339 DIN3 GVSS 0 nch W=0.84U L=0.24U
M8 GVSS DIN4 N1N339 0 nch W=0.84U L=0.24U
M5 N1N339 DIN1 Q 0 nch W=0.84U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai13s3 Q DIN1 DIN2 DIN3 DIN4
M1 N1N330 DIN2 VDD VDD pch W=1.8U L=0.24U
M6 N1N339 DIN2 GVSS 0 nch W=0.9U L=0.24U
M2 N1N332 DIN3 N1N330 VDD pch W=1.8U L=0.24U
M3 N1N334 DIN4 N1N332 VDD pch W=1.8U L=0.24U
M4 VDD DIN1 N1N334 VDD pch W=0.66U L=0.24U
M7 N1N339 DIN3 GVSS 0 nch W=0.9U L=0.24U
M8 GVSS DIN4 N1N339 0 nch W=0.9U L=0.24U
M5 N1N339 DIN1 N1N334 0 nch W=0.9U L=0.24U
M10 N1N383 N1N334 GVSS 0 nch W=1.2U L=0.24U
M12 Q N1N383 GVSS 0 nch W=2U L=0.24U
M9 N1N383 N1N334 VDD VDD pch W=2.3U L=0.24U
M11 Q N1N383 VDD VDD pch W=4.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai211s1 Q DIN1 DIN2 DIN3 DIN4
M6 N1N469 DIN3 N1N444 0 nch W=0.8U L=0.24U
M1 N1N435 DIN1 VDD VDD pch W=1.8U L=0.24U
M2 Q DIN2 N1N435 VDD pch W=1.8U L=0.24U
M3 Q DIN3 VDD VDD pch W=0.7U L=0.24U
M4 VDD DIN4 Q VDD pch W=0.7U L=0.24U
M7 N1N444 DIN1 GVSS 0 nch W=0.8U L=0.24U
M5 N1N469 DIN4 Q 0 nch W=0.7U L=0.24U
M8 GVSS DIN2 N1N444 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai211s2 Q DIN1 DIN2 DIN3 DIN4
M6 N1N469 DIN3 N1N444 0 nch W=1.2U L=0.24U
M1 N1N435 DIN1 VDD VDD pch W=2.9U L=0.24U
M2 Q DIN2 N1N435 VDD pch W=2.8U L=0.24U
M3 Q DIN3 VDD VDD pch W=1.1U L=0.24U
M4 VDD DIN4 Q VDD pch W=1.1U L=0.24U
M7 N1N444 DIN1 GVSS 0 nch W=1.3U L=0.24U
M5 N1N469 DIN4 Q 0 nch W=1.1U L=0.24U
M8 GVSS DIN2 N1N444 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai211s3 Q DIN1 DIN2 DIN3 DIN4
M6 N1N326 DIN3 N1N327 0 nch W=0.9U L=0.24U
M1 N1N332 DIN1 VDD VDD pch W=2U L=0.24U
M2 N1N329 DIN2 N1N332 VDD pch W=2U L=0.24U
M3 N1N329 DIN3 VDD VDD pch W=0.8U L=0.24U
M4 VDD DIN4 N1N329 VDD pch W=0.8U L=0.24U
M7 N1N327 DIN1 GVSS 0 nch W=0.9U L=0.24U
M5 N1N326 DIN4 N1N329 0 nch W=0.8U L=0.24U
M8 GVSS DIN2 N1N327 0 nch W=0.9U L=0.24U
M10 N1N374 N1N329 GVSS 0 nch W=1.2U L=0.24U
M9 N1N374 N1N329 VDD VDD pch W=2U L=0.24U
M11 Q N1N374 VDD VDD pch W=4.3U L=0.24U
M12 Q N1N374 GVSS 0 nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai21s1 Q DIN1 DIN2 DIN3
M5 N1N261 DIN2 GVSS 0 nch W=0.6U L=0.24U
M1 Q DIN3 VDD VDD pch W=0.7U L=0.24U
M2 VDD DIN1 N1N257 VDD pch W=1.7U L=0.24U
M3 N1N257 DIN2 Q VDD pch W=1.7U L=0.24U
M4 Q DIN3 N1N261 0 nch W=0.6U L=0.24U
M6 GVSS DIN1 N1N261 0 nch W=0.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai21s2 Q DIN1 DIN2 DIN3
M5 N1N284 DIN2 GVSS 0 nch W=1U L=0.24U
M1 Q DIN3 VDD VDD pch W=1.2U L=0.24U
M2 VDD DIN1 N1N257 VDD pch W=2.8U L=0.24U
M3 N1N257 DIN2 Q VDD pch W=2.7U L=0.24U
M4 Q DIN3 N1N284 0 nch W=1U L=0.24U
M6 GVSS DIN1 N1N284 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai21s3 Q DIN1 DIN2 DIN3
M5 N1N284 DIN2 GVSS 0 nch W=2U L=0.24U
M1 Q DIN3 VDD VDD pch W=2.1U L=0.24U
M2 VDD DIN1 N1N257 VDD pch W=5.6U L=0.24U
M3 N1N257 DIN2 Q VDD pch W=5.4U L=0.24U
M4 Q DIN3 N1N284 0 nch W=2U L=0.24U
M6 GVSS DIN1 N1N284 0 nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai221s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M7 N1N283 DIN3 N1N292 0 nch W=0.8U L=0.24U
M1 N1N263 DIN1 VDD VDD pch W=1.8U L=0.24U
M2 Q DIN2 N1N263 VDD pch W=1.8U L=0.24U
M3 VDD DIN3 N1N290 VDD pch W=1.8U L=0.24U
M5 VDD DIN5 Q VDD pch W=0.8U L=0.24U
M4 N1N290 DIN4 Q VDD pch W=1.8U L=0.24U
M9 N1N292 DIN1 GVSS 0 nch W=0.8U L=0.24U
M10 GVSS DIN2 N1N292 0 nch W=0.8U L=0.24U
M8 N1N292 DIN4 N1N283 0 nch W=0.8U L=0.24U
M6 N1N283 DIN5 Q 0 nch W=0.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai221s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M7 N1N283 DIN3 N1N292 0 nch W=1.2U L=0.24U
M1 N1N263 DIN1 VDD VDD pch W=2.9U L=0.24U
M2 Q DIN2 N1N263 VDD pch W=2.8U L=0.24U
M3 VDD DIN3 N1N290 VDD pch W=2.9U L=0.24U
M5 VDD DIN5 Q VDD pch W=1.1U L=0.24U
M4 N1N290 DIN4 Q VDD pch W=2.8U L=0.24U
M9 N1N292 DIN1 GVSS 0 nch W=1.3U L=0.24U
M10 GVSS DIN2 N1N292 0 nch W=1.3U L=0.24U
M8 N1N292 DIN4 N1N283 0 nch W=1.2U L=0.24U
M6 N1N283 DIN5 Q 0 nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai221s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M7 N1N283 DIN3 N1N292 0 nch W=0.9U L=0.24U
M1 N1N263 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N265 DIN2 N1N263 VDD pch W=2U L=0.24U
M3 VDD DIN3 N1N290 VDD pch W=2.1U L=0.24U
M5 VDD DIN5 N1N265 VDD pch W=0.8U L=0.24U
M4 N1N290 DIN4 N1N265 VDD pch W=2U L=0.24U
M9 N1N292 DIN1 GVSS 0 nch W=1U L=0.24U
M10 GVSS DIN2 N1N292 0 nch W=1U L=0.24U
M8 N1N292 DIN4 N1N283 0 nch W=0.9U L=0.24U
M6 N1N283 DIN5 N1N265 0 nch W=0.8U L=0.24U
M12 N1N351 N1N265 GVSS 0 nch W=1.3U L=0.24U
M11 N1N351 N1N265 VDD VDD pch W=2.2U L=0.24U
M13 Q N1N351 VDD VDD pch W=4.5U L=0.24U
M14 Q N1N351 GVSS 0 nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai2222s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8
M3 N1N271 DIN2 N1N273 0 nch W=0.7U L=0.24U
M6 N1N271 DIN1 N1N276 VDD pch W=1U L=0.24U
M2 N1N271 DIN3 N1N269 VDD pch W=1U L=0.24U
M4 N1N273 DIN3 GVSS 0 nch W=0.7U L=0.24U
M1 N1N269 DIN4 VDD VDD pch W=1U L=0.24U
M5 N1N276 DIN2 VDD VDD pch W=1U L=0.24U
M7 N1N271 DIN1 N1N273 0 nch W=0.7U L=0.24U
M8 N1N273 DIN4 GVSS 0 nch W=0.7U L=0.24U
M11 N1N315 DIN6 N1N319 0 nch W=0.7U L=0.24U
M9 N1N354 DIN8 VDD VDD pch W=1U L=0.24U
M10 N1N315 DIN7 N1N354 VDD pch W=1U L=0.24U
M12 N1N319 DIN7 GVSS 0 nch W=0.7U L=0.24U
M16 N1N319 DIN8 GVSS 0 nch W=0.7U L=0.24U
M15 N1N315 DIN5 N1N319 0 nch W=0.7U L=0.24U
M13 N1N325 DIN6 VDD VDD pch W=1U L=0.24U
M14 N1N315 DIN5 N1N325 VDD pch W=1U L=0.24U
M19 N1N328 N1N271 GVSS 0 nch W=0.6U L=0.24U
M18 N1N328 N1N271 N1N357 VDD pch W=1.5U L=0.24U
M17 VDD N1N315 N1N357 VDD pch W=1.5U L=0.24U
M20 N1N328 N1N315 GVSS 0 nch W=0.6U L=0.24U
M22 Q N1N328 GVSS 0 nch W=1U L=0.24U
M21 Q N1N328 VDD VDD pch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai2222s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8
M3 N1N271 DIN2 N1N273 0 nch W=0.7U L=0.24U
M6 N1N271 DIN1 N1N276 VDD pch W=1U L=0.24U
M2 N1N271 DIN3 N1N269 VDD pch W=1U L=0.24U
M4 N1N273 DIN3 GVSS 0 nch W=0.7U L=0.24U
M1 N1N269 DIN4 VDD VDD pch W=1U L=0.24U
M5 N1N276 DIN2 VDD VDD pch W=1U L=0.24U
M7 N1N271 DIN1 N1N273 0 nch W=0.7U L=0.24U
M8 N1N273 DIN4 GVSS 0 nch W=0.7U L=0.24U
M11 N1N315 DIN6 N1N319 0 nch W=0.7U L=0.24U
M9 N1N354 DIN8 VDD VDD pch W=1U L=0.24U
M10 N1N315 DIN7 N1N354 VDD pch W=1U L=0.24U
M12 N1N319 DIN7 GVSS 0 nch W=0.7U L=0.24U
M16 N1N319 DIN8 GVSS 0 nch W=0.7U L=0.24U
M15 N1N315 DIN5 N1N319 0 nch W=0.7U L=0.24U
M13 N1N325 DIN6 VDD VDD pch W=1U L=0.24U
M14 N1N315 DIN5 N1N325 VDD pch W=1U L=0.24U
M19 N1N328 N1N271 GVSS 0 nch W=0.9U L=0.24U
M18 N1N328 N1N271 N1N357 VDD pch W=2.2U L=0.24U
M17 VDD N1N315 N1N357 VDD pch W=2.2U L=0.24U
M20 N1N328 N1N315 GVSS 0 nch W=0.9U L=0.24U
M22 Q N1N328 GVSS 0 nch W=1.4U L=0.24U
M21 Q N1N328 VDD VDD pch W=3.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai2222s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8
M3 N1N271 DIN2 N1N273 0 nch W=1.4U L=0.24U
M6 N1N271 DIN1 N1N276 VDD pch W=2U L=0.24U
M2 N1N271 DIN3 N1N269 VDD pch W=2U L=0.24U
M4 N1N273 DIN3 GVSS 0 nch W=1.4U L=0.24U
M1 N1N269 DIN4 VDD VDD pch W=2U L=0.24U
M5 N1N276 DIN2 VDD VDD pch W=2U L=0.24U
M7 N1N271 DIN1 N1N273 0 nch W=1.4U L=0.24U
M8 N1N273 DIN4 GVSS 0 nch W=1.4U L=0.24U
M11 N1N315 DIN6 N1N319 0 nch W=1.4U L=0.24U
M9 N1N354 DIN8 VDD VDD pch W=2U L=0.24U
M10 N1N315 DIN7 N1N354 VDD pch W=2U L=0.24U
M12 N1N319 DIN7 GVSS 0 nch W=1.4U L=0.24U
M16 N1N319 DIN8 GVSS 0 nch W=1.4U L=0.24U
M15 N1N315 DIN5 N1N319 0 nch W=1.4U L=0.24U
M13 N1N325 DIN6 VDD VDD pch W=2U L=0.24U
M14 N1N315 DIN5 N1N325 VDD pch W=2U L=0.24U
M19 N1N328 N1N271 GVSS 0 nch W=1.5U L=0.24U
M18 N1N328 N1N271 N1N357 VDD pch W=3.4U L=0.24U
M17 VDD N1N315 N1N357 VDD pch W=3.4U L=0.24U
M20 N1N328 N1N315 GVSS 0 nch W=1.5U L=0.24U
M22 Q N1N328 GVSS 0 nch W=2.1U L=0.24U
M21 Q N1N328 VDD VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai222s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN5 N1N334 0 nch W=0.9U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=1.9U L=0.24U
M4 Q DIN2 N1N323 VDD pch W=1.9U L=0.24U
M2 VDD DIN3 N1N325 VDD pch W=1.9U L=0.24U
M5 N1N325 DIN4 Q VDD pch W=1.9U L=0.24U
M3 VDD DIN5 N1N327 VDD pch W=1.9U L=0.24U
M6 N1N327 DIN6 Q VDD pch W=1.9U L=0.24U
M9 N1N334 DIN3 N1N338 0 nch W=0.9U L=0.24U
M11 N1N338 DIN1 GVSS 0 nch W=0.9U L=0.24U
M12 GVSS DIN2 N1N338 0 nch W=0.9U L=0.24U
M10 N1N338 DIN4 N1N334 0 nch W=0.9U L=0.24U
M8 N1N334 DIN6 Q 0 nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai222s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N329 DIN5 N1N334 0 nch W=0.9U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=2U L=0.24U
M4 N1N329 DIN2 N1N323 VDD pch W=1.9U L=0.24U
M2 VDD DIN3 N1N325 VDD pch W=2U L=0.24U
M5 N1N325 DIN4 N1N329 VDD pch W=1.9U L=0.24U
M3 VDD DIN5 N1N327 VDD pch W=2U L=0.24U
M6 N1N327 DIN6 N1N329 VDD pch W=1.9U L=0.24U
M9 N1N334 DIN3 N1N338 0 nch W=0.9U L=0.24U
M11 N1N338 DIN1 GVSS 0 nch W=1U L=0.24U
M12 GVSS DIN2 N1N338 0 nch W=1U L=0.24U
M10 N1N338 DIN4 N1N334 0 nch W=0.9U L=0.24U
M8 N1N334 DIN6 N1N329 0 nch W=0.9U L=0.24U
M14 N1N370 N1N329 GVSS 0 nch W=0.6U L=0.24U
M13 N1N370 N1N329 VDD VDD pch W=1.3U L=0.24U
M15 Q N1N370 VDD VDD pch W=2.4U L=0.24U
M16 Q N1N370 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai222s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N329 DIN5 N1N334 0 nch W=0.9U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=2.04U L=0.24U
M4 N1N329 DIN2 N1N323 VDD pch W=1.9U L=0.24U
M2 VDD DIN3 N1N325 VDD pch W=2.04U L=0.24U
M5 N1N325 DIN4 N1N329 VDD pch W=1.9U L=0.24U
M3 VDD DIN5 N1N327 VDD pch W=2.04U L=0.24U
M6 N1N327 DIN6 N1N329 VDD pch W=1.9U L=0.24U
M9 N1N334 DIN3 N1N338 0 nch W=1U L=0.24U
M11 N1N338 DIN1 GVSS 0 nch W=1.1U L=0.24U
M12 GVSS DIN2 N1N338 0 nch W=1.1U L=0.24U
M10 N1N338 DIN4 N1N334 0 nch W=1U L=0.24U
M8 N1N334 DIN6 N1N329 0 nch W=0.9U L=0.24U
M14 N1N372 N1N329 GVSS 0 nch W=1U L=0.24U
M13 N1N372 N1N329 VDD VDD pch W=2.2U L=0.24U
M16 Q N1N372 GVSS 0 nch W=2.1U L=0.24U
M15 Q N1N372 VDD VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai22s1 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N278 0 nch W=0.64U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=1.7U L=0.24U
M2 Q DIN2 N1N258 VDD pch W=1.7U L=0.24U
M4 N1N260 DIN4 Q VDD pch W=1.7U L=0.24U
M3 VDD DIN3 N1N260 VDD pch W=1.7U L=0.24U
M6 N1N278 DIN3 GVSS 0 nch W=0.64U L=0.24U
M8 GVSS DIN4 N1N278 0 nch W=0.64U L=0.24U
M7 N1N278 DIN2 Q 0 nch W=0.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai22s2 Q DIN1 DIN2 DIN3 DIN4
M5 Q DIN1 N1N278 0 nch W=1.02U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=2.6U L=0.24U
M2 Q DIN2 N1N258 VDD pch W=2.6U L=0.24U
M4 N1N260 DIN4 Q VDD pch W=2.6U L=0.24U
M3 VDD DIN3 N1N260 VDD pch W=2.6U L=0.24U
M6 N1N278 DIN3 GVSS 0 nch W=1.02U L=0.24U
M8 GVSS DIN4 N1N278 0 nch W=1.02U L=0.24U
M7 N1N278 DIN2 Q 0 nch W=1.02U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai22s3 Q DIN1 DIN2 DIN3 DIN4
M5 N1N268 DIN1 N1N278 0 nch W=0.8U L=0.24U
M1 N1N258 DIN1 VDD VDD pch W=1.8U L=0.24U
M2 N1N268 DIN2 N1N258 VDD pch W=1.7U L=0.24U
M4 N1N260 DIN4 N1N268 VDD pch W=1.7U L=0.24U
M3 VDD DIN3 N1N260 VDD pch W=1.8U L=0.24U
M6 N1N278 DIN3 GVSS 0 nch W=0.8U L=0.24U
M8 GVSS DIN4 N1N278 0 nch W=0.8U L=0.24U
M7 N1N278 DIN2 N1N268 0 nch W=0.8U L=0.24U
M10 N1N295 N1N268 GVSS 0 nch W=1.2U L=0.24U
M9 N1N295 N1N268 VDD VDD pch W=2.3U L=0.24U
M11 Q N1N295 VDD VDD pch W=4.3U L=0.24U
M12 Q N1N295 GVSS 0 nch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai24s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N311 0 nch W=0.8U L=0.24U
M1 N1N301 DIN1 VDD VDD pch W=2.3U L=0.24U
M3 Q DIN2 N1N301 VDD pch W=2.1U L=0.24U
M2 VDD DIN3 N1N303 VDD pch W=4.4U L=0.24U
M4 N1N303 DIN4 N1N305 VDD pch W=4.4U L=0.24U
M5 N1N305 DIN5 N1N307 VDD pch W=4.2U L=0.24U
M6 N1N307 DIN6 Q VDD pch W=4.2U L=0.24U
M9 N1N311 DIN3 GVSS 0 nch W=0.8U L=0.24U
M8 N1N311 DIN2 Q 0 nch W=0.8U L=0.24U
M10 GVSS DIN6 N1N311 0 nch W=0.8U L=0.24U
M11 N1N311 DIN4 GVSS 0 nch W=0.8U L=0.24U
M12 GVSS DIN5 N1N311 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai24s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N311 0 nch W=1.3U L=0.24U
M1 N1N301 DIN1 VDD VDD pch W=3.5U L=0.24U
M3 Q DIN2 N1N301 VDD pch W=3.4U L=0.24U
M2 VDD DIN3 N1N303 VDD pch W=6.6U L=0.24U
M4 N1N303 DIN4 N1N305 VDD pch W=6.6U L=0.24U
M5 N1N305 DIN5 N1N307 VDD pch W=6.4U L=0.24U
M6 N1N307 DIN6 Q VDD pch W=6.4U L=0.24U
M9 N1N311 DIN3 GVSS 0 nch W=1.3U L=0.24U
M8 N1N311 DIN2 Q 0 nch W=1.3U L=0.24U
M10 GVSS DIN6 N1N311 0 nch W=1.3U L=0.24U
M11 N1N311 DIN4 GVSS 0 nch W=1.3U L=0.24U
M12 GVSS DIN5 N1N311 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai24s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N311 0 nch W=2.14U L=0.24U
M1 N1N301 DIN1 VDD VDD pch W=5.3U L=0.24U
M3 Q DIN2 N1N301 VDD pch W=5.2U L=0.24U
M2 VDD DIN3 N1N303 VDD pch W=9.9U L=0.24U
M4 N1N303 DIN4 N1N305 VDD pch W=9.9U L=0.24U
M5 N1N305 DIN5 N1N307 VDD pch W=9.8U L=0.24U
M6 N1N307 DIN6 Q VDD pch W=9.8U L=0.24U
M9 N1N311 DIN3 GVSS 0 nch W=2.14U L=0.24U
M8 N1N311 DIN2 Q 0 nch W=2.14U L=0.24U
M10 GVSS DIN6 N1N311 0 nch W=2.14U L=0.24U
M11 N1N311 DIN4 GVSS 0 nch W=2.14U L=0.24U
M12 GVSS DIN5 N1N311 0 nch W=2.14U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai321s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M12 N1N284 DIN3 GVSS 0 nch W=1.1U L=0.24U
M6 Q DIN3 N1N257 VDD pch W=2.9U L=0.24U
M5 N1N257 DIN2 N1N256 VDD pch W=3U L=0.24U
M4 N1N256 DIN1 VDD VDD pch W=3.1U L=0.24U
M3 Q DIN6 VDD VDD pch W=1U L=0.24U
M2 Q DIN5 N1N278 VDD pch W=2U L=0.24U
M11 N1N284 DIN1 GVSS 0 nch W=1.1U L=0.24U
M9 N1N282 DIN4 N1N284 0 nch W=1U L=0.24U
M10 N1N284 DIN2 GVSS 0 nch W=1.1U L=0.24U
M7 Q DIN6 N1N282 0 nch W=1U L=0.24U
M8 N1N282 DIN5 N1N284 0 nch W=1U L=0.24U
M1 N1N278 DIN4 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai321s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M12 N1N284 DIN3 GVSS 0 nch W=1.1U L=0.24U
M6 N1N280 DIN3 N1N257 VDD pch W=2.9U L=0.24U
M5 N1N257 DIN2 N1N256 VDD pch W=3U L=0.24U
M4 N1N256 DIN1 VDD VDD pch W=3.1U L=0.24U
M3 N1N280 DIN6 VDD VDD pch W=1U L=0.24U
M2 N1N280 DIN5 N1N278 VDD pch W=2U L=0.24U
M1 N1N278 DIN4 VDD VDD pch W=2U L=0.24U
M11 N1N284 DIN1 GVSS 0 nch W=1.1U L=0.24U
M9 N1N282 DIN4 N1N284 0 nch W=1U L=0.24U
M10 N1N284 DIN2 GVSS 0 nch W=1.1U L=0.24U
M7 N1N280 DIN6 N1N282 0 nch W=1U L=0.24U
M8 N1N282 DIN5 N1N284 0 nch W=1U L=0.24U
M14 N1N325 N1N280 GVSS 0 nch W=0.64U L=0.24U
M13 N1N325 N1N280 VDD VDD pch W=1.4U L=0.24U
M15 Q N1N325 VDD VDD pch W=2.4U L=0.24U
M16 Q N1N325 GVSS 0 nch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai321s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M12 N1N284 DIN3 GVSS 0 nch W=1.2U L=0.24U
M6 N1N280 DIN3 N1N257 VDD pch W=2.9U L=0.24U
M5 N1N257 DIN2 N1N256 VDD pch W=3U L=0.24U
M4 N1N256 DIN1 VDD VDD pch W=3.1U L=0.24U
M3 N1N280 DIN6 VDD VDD pch W=1U L=0.24U
M2 N1N280 DIN5 N1N278 VDD pch W=2U L=0.24U
M1 N1N278 DIN4 VDD VDD pch W=2U L=0.24U
M11 N1N284 DIN1 GVSS 0 nch W=1.2U L=0.24U
M9 N1N282 DIN4 N1N284 0 nch W=1.1U L=0.24U
M10 N1N284 DIN2 GVSS 0 nch W=1.2U L=0.24U
M7 N1N280 DIN6 N1N282 0 nch W=1U L=0.24U
M8 N1N282 DIN5 N1N284 0 nch W=1.1U L=0.24U
M14 N1N322 N1N280 GVSS 0 nch W=1.1U L=0.24U
M13 N1N322 N1N280 VDD VDD pch W=2.52U L=0.24U
M15 Q N1N322 VDD VDD pch W=4.2U L=0.24U
M16 Q N1N322 GVSS 0 nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai322s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M3 Q DIN6 N1N322 0 nch W=1U L=0.24U
M1 N1N307 DIN4 VDD VDD pch W=1.5U L=0.24U
M2 Q DIN5 N1N307 VDD pch W=1.5U L=0.24U
M6 N1N311 DIN6 VDD VDD pch W=1.5U L=0.24U
M7 Q DIN7 N1N311 VDD pch W=1.5U L=0.24U
M4 N1N322 DIN5 N1N326 0 nch W=1U L=0.24U
M5 N1N326 DIN2 GVSS 0 nch W=1U L=0.24U
M8 Q DIN7 N1N322 0 nch W=1U L=0.24U
M9 N1N322 DIN4 N1N326 0 nch W=1U L=0.24U
M10 N1N326 DIN1 GVSS 0 nch W=1U L=0.24U
M11 N1N318 DIN1 VDD VDD pch W=2.3U L=0.24U
M12 N1N320 DIN2 N1N318 VDD pch W=2.3U L=0.24U
M13 Q DIN3 N1N320 VDD pch W=2.3U L=0.24U
M14 N1N326 DIN3 GVSS 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai322s2 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M3 N1N309 DIN6 N1N322 0 nch W=1U L=0.24U
M1 N1N307 DIN4 VDD VDD pch W=1.5U L=0.24U
M2 N1N309 DIN5 N1N307 VDD pch W=1.5U L=0.24U
M6 N1N311 DIN6 VDD VDD pch W=1.5U L=0.24U
M7 N1N309 DIN7 N1N311 VDD pch W=1.5U L=0.24U
M4 N1N322 DIN5 N1N326 0 nch W=1.1U L=0.24U
M5 N1N326 DIN2 GVSS 0 nch W=1.1U L=0.24U
M8 N1N309 DIN7 N1N322 0 nch W=1U L=0.24U
M9 N1N322 DIN4 N1N326 0 nch W=1.1U L=0.24U
M10 N1N326 DIN1 GVSS 0 nch W=1.1U L=0.24U
M11 N1N318 DIN1 VDD VDD pch W=2.3U L=0.24U
M12 N1N320 DIN2 N1N318 VDD pch W=2.3U L=0.24U
M13 N1N309 DIN3 N1N320 VDD pch W=2.3U L=0.24U
M14 N1N326 DIN3 GVSS 0 nch W=1.1U L=0.24U
M15 N1N360 N1N309 VDD VDD pch W=2.7U L=0.24U
M16 N1N360 N1N309 GVSS 0 nch W=1.1U L=0.24U
M18 Q N1N360 GVSS 0 nch W=2.3U L=0.24U
M17 Q N1N360 VDD VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai322s3 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 Q
M3 N1N309 DIN6 N1N322 0 nch W=1.1U L=0.24U
M1 N1N307 DIN4 VDD VDD pch W=1.8U L=0.24U
M2 N1N309 DIN5 N1N307 VDD pch W=1.8U L=0.24U
M6 N1N311 DIN6 VDD VDD pch W=1.8U L=0.24U
M7 N1N309 DIN7 N1N311 VDD pch W=1.8U L=0.24U
M4 N1N322 DIN5 N1N326 0 nch W=1.3U L=0.24U
M5 N1N326 DIN2 GVSS 0 nch W=1.3U L=0.24U
M8 N1N309 DIN7 N1N322 0 nch W=1.1U L=0.24U
M9 N1N322 DIN4 N1N326 0 nch W=1.3U L=0.24U
M10 N1N326 DIN1 GVSS 0 nch W=1.3U L=0.24U
M11 N1N318 DIN1 VDD VDD pch W=2.7U L=0.24U
M12 N1N320 DIN2 N1N318 VDD pch W=2.7U L=0.24U
M13 N1N309 DIN3 N1N320 VDD pch W=2.7U L=0.24U
M14 N1N326 DIN3 GVSS 0 nch W=1.3U L=0.24U
M15 N1N360 N1N309 VDD VDD pch W=4.2U L=0.24U
M16 N1N360 N1N309 GVSS 0 nch W=1.7U L=0.24U
M18 Q N1N360 GVSS 0 nch W=3.6U L=0.24U
M17 Q N1N360 VDD VDD pch W=6.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai32s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN5 N1N333 0 nch W=0.8U L=0.24U
M1 N1N321 DIN1 VDD VDD pch W=3.2U L=0.24U
M2 N1N323 DIN2 N1N321 VDD pch W=3.2U L=0.24U
M3 Q DIN3 N1N323 VDD pch W=3.2U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2.1U L=0.24U
M5 N1N327 DIN5 Q VDD pch W=2.1U L=0.24U
M8 N1N333 DIN1 GVSS 0 nch W=0.8U L=0.24U
M9 GVSS DIN2 N1N333 0 nch W=0.8U L=0.24U
M7 N1N333 DIN4 Q 0 nch W=0.8U L=0.24U
M10 GVSS DIN3 N1N333 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai32s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 Q DIN5 N1N333 0 nch W=1U L=0.24U
M1 N1N321 DIN1 VDD VDD pch W=4.1U L=0.24U
M2 N1N323 DIN2 N1N321 VDD pch W=4U L=0.24U
M3 Q DIN3 N1N323 VDD pch W=3.9U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2.6U L=0.24U
M5 N1N327 DIN5 Q VDD pch W=2.5U L=0.24U
M8 N1N333 DIN1 GVSS 0 nch W=1U L=0.24U
M9 GVSS DIN2 N1N333 0 nch W=1U L=0.24U
M7 N1N333 DIN4 Q 0 nch W=1U L=0.24U
M10 GVSS DIN3 N1N333 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai32s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M6 N1N325 DIN5 N1N333 0 nch W=0.9U L=0.24U
M1 N1N321 DIN1 VDD VDD pch W=3.1U L=0.24U
M2 N1N323 DIN2 N1N321 VDD pch W=3.1U L=0.24U
M3 N1N325 DIN3 N1N323 VDD pch W=3.1U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2U L=0.24U
M5 N1N327 DIN5 N1N325 VDD pch W=2U L=0.24U
M8 N1N333 DIN1 GVSS 0 nch W=0.9U L=0.24U
M9 GVSS DIN2 N1N333 0 nch W=0.9U L=0.24U
M7 N1N333 DIN4 N1N325 0 nch W=0.9U L=0.24U
M10 GVSS DIN3 N1N333 0 nch W=0.9U L=0.24U
M11 N1N369 N1N325 VDD VDD pch W=2.5U L=0.24U
M13 Q N1N369 VDD VDD pch W=4.5U L=0.24U
M12 N1N369 N1N325 GVSS 0 nch W=1.4U L=0.24U
M14 Q N1N369 GVSS 0 nch W=2.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai33s1 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 Q DIN1 N1N335 0 nch W=0.9U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=3.1U L=0.24U
M2 N1N331 DIN2 N1N323 VDD pch W=3U L=0.24U
M3 Q DIN3 N1N331 VDD pch W=2.9U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=3.1U L=0.24U
M5 N1N327 DIN5 N1N329 VDD pch W=3U L=0.24U
M6 N1N329 DIN6 Q VDD pch W=2.9U L=0.24U
M8 N1N335 DIN4 GVSS 0 nch W=1.1U L=0.24U
M9 Q DIN2 N1N335 0 nch W=0.9U L=0.24U
M10 N1N335 DIN5 GVSS 0 nch W=1.1U L=0.24U
M11 N1N335 DIN3 Q 0 nch W=0.9U L=0.24U
M12 GVSS DIN6 N1N335 0 nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai33s2 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N333 DIN1 N1N335 0 nch W=0.8U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N331 DIN2 N1N323 VDD pch W=1.9U L=0.24U
M3 N1N333 DIN3 N1N331 VDD pch W=1.9U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2.1U L=0.24U
M5 N1N327 DIN5 N1N329 VDD pch W=1.9U L=0.24U
M6 N1N329 DIN6 N1N333 VDD pch W=1.9U L=0.24U
M8 N1N335 DIN4 GVSS 0 nch W=0.9U L=0.24U
M9 N1N333 DIN2 N1N335 0 nch W=0.8U L=0.24U
M10 N1N335 DIN5 GVSS 0 nch W=0.9U L=0.24U
M11 N1N335 DIN3 N1N333 0 nch W=0.8U L=0.24U
M12 GVSS DIN6 N1N335 0 nch W=0.9U L=0.24U
M13 N1N383 N1N333 VDD VDD pch W=1.1U L=0.24U
M14 N1N383 N1N333 GVSS 0 nch W=0.6U L=0.24U
M15 Q N1N383 VDD VDD pch W=2.4U L=0.24U
M16 Q N1N383 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_oai33s3 Q DIN1 DIN2 DIN3 DIN4 DIN5 DIN6
M7 N1N333 DIN1 N1N335 0 nch W=0.8U L=0.24U
M1 N1N323 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N331 DIN2 N1N323 VDD pch W=1.9U L=0.24U
M3 N1N333 DIN3 N1N331 VDD pch W=1.9U L=0.24U
M4 VDD DIN4 N1N327 VDD pch W=2.1U L=0.24U
M5 N1N327 DIN5 N1N329 VDD pch W=1.9U L=0.24U
M6 N1N329 DIN6 N1N333 VDD pch W=1.9U L=0.24U
M8 N1N335 DIN4 GVSS 0 nch W=0.9U L=0.24U
M9 N1N333 DIN2 N1N335 0 nch W=0.8U L=0.24U
M10 N1N335 DIN5 GVSS 0 nch W=0.9U L=0.24U
M11 N1N335 DIN3 N1N333 0 nch W=0.8U L=0.24U
M12 GVSS DIN6 N1N335 0 nch W=0.9U L=0.24U
M13 N1N383 N1N333 VDD VDD pch W=2U L=0.24U
M14 N1N383 N1N333 GVSS 0 nch W=1U L=0.24U
M15 Q N1N383 VDD VDD pch W=4.2U L=0.24U
M16 Q N1N383 GVSS 0 nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or2s1 Q DIN1 DIN2
M3 N1N441 DIN1 GVSS 0 nch W=0.7U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=1.6U L=0.24U
M2 N1N441 DIN2 N1N428 VDD pch W=1.6U L=0.24U
M4 N1N441 DIN2 GVSS 0 nch W=0.7U L=0.24U
M6 Q N1N441 GVSS 0 nch W=1.3U L=0.24U
M5 Q N1N441 VDD VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or2s2 Q DIN1 DIN2
M3 N1N441 DIN1 GVSS 0 nch W=1.1U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=3U L=0.24U
M2 N1N441 DIN2 N1N428 VDD pch W=3U L=0.24U
M4 N1N441 DIN2 GVSS 0 nch W=1.1U L=0.24U
M6 Q N1N441 GVSS 0 nch W=3.5U L=0.24U
M5 Q N1N441 VDD VDD pch W=4.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or2s3 Q DIN1 DIN2
M3 N1N441 DIN1 GVSS 0 nch W=2.2U L=0.24U
M1 N1N428 DIN1 VDD VDD pch W=5.8U L=0.24U
M2 N1N441 DIN2 N1N428 VDD pch W=5.8U L=0.24U
M4 N1N441 DIN2 GVSS 0 nch W=2.2U L=0.24U
M6 Q N1N441 GVSS 0 nch W=6.2U L=0.24U
M5 Q N1N441 VDD VDD pch W=7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or3s1 Q DIN1 DIN2 DIN3
M4 N1N434 DIN1 GVSS 0 nch W=0.7U L=0.24U
M1 N1N430 DIN1 VDD VDD pch W=3.16U L=0.24U
M2 N1N432 DIN2 N1N430 VDD pch W=3.16U L=0.24U
M3 N1N434 DIN3 N1N432 VDD pch W=3.16U L=0.24U
M5 N1N434 DIN2 GVSS 0 nch W=0.7U L=0.24U
M6 N1N434 DIN3 GVSS 0 nch W=0.7U L=0.24U
M7 Q N1N434 VDD VDD pch W=2.1U L=0.24U
M8 Q N1N434 GVSS 0 nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or3s2 Q DIN1 DIN2 DIN3
M4 N1N434 DIN1 GVSS 0 nch W=1.1U L=0.24U
M1 N1N430 DIN1 VDD VDD pch W=4.2U L=0.24U
M2 N1N432 DIN2 N1N430 VDD pch W=4.1U L=0.24U
M3 N1N434 DIN3 N1N432 VDD pch W=4U L=0.24U
M5 N1N434 DIN2 GVSS 0 nch W=1.1U L=0.24U
M6 N1N434 DIN3 GVSS 0 nch W=1.1U L=0.24U
M7 Q N1N434 VDD VDD pch W=5.2U L=0.24U
M8 Q N1N434 GVSS 0 nch W=4.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or3s3 Q DIN1 DIN2 DIN3
M4 N1N434 DIN1 GVSS 0 nch W=2U L=0.24U
M1 N1N430 DIN1 VDD VDD pch W=8.5U L=0.24U
M2 N1N432 DIN2 N1N430 VDD pch W=7.8U L=0.24U
M3 N1N434 DIN3 N1N432 VDD pch W=6.2U L=0.24U
M5 N1N434 DIN2 GVSS 0 nch W=2U L=0.24U
M6 N1N434 DIN3 GVSS 0 nch W=2U L=0.24U
M7 Q N1N434 VDD VDD pch W=7.1U L=0.24U
M8 Q N1N434 GVSS 0 nch W=6.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or4s1 Q DIN1 DIN2 DIN3 DIN4
M5 N1N438 DIN1 GVSS 0 nch W=0.7U L=0.24U
M1 N1N432 DIN1 VDD VDD pch W=4.5U L=0.24U
M2 N1N434 DIN2 N1N432 VDD pch W=4.2U L=0.24U
M3 N1N436 DIN3 N1N434 VDD pch W=4.1U L=0.24U
M4 N1N438 DIN4 N1N436 VDD pch W=3.1U L=0.24U
M6 N1N438 DIN2 GVSS 0 nch W=0.7U L=0.24U
M7 N1N438 DIN3 GVSS 0 nch W=0.7U L=0.24U
M8 N1N438 DIN4 GVSS 0 nch W=0.7U L=0.24U
M9 Q N1N438 VDD VDD pch W=2.3U L=0.24U
M10 Q N1N438 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or4s2 Q DIN1 DIN2 DIN3 DIN4
M5 N1N438 DIN1 GVSS 0 nch W=1.56U L=0.24U
M1 N1N432 DIN1 VDD VDD pch W=9.5U L=0.24U
M2 N1N434 DIN2 N1N432 VDD pch W=9.2U L=0.24U
M3 N1N436 DIN3 N1N434 VDD pch W=9U L=0.24U
M4 N1N438 DIN4 N1N436 VDD pch W=8.5U L=0.24U
M6 N1N438 DIN2 GVSS 0 nch W=1.56U L=0.24U
M7 N1N438 DIN3 GVSS 0 nch W=1.56U L=0.24U
M8 N1N438 DIN4 GVSS 0 nch W=1.56U L=0.24U
M9 Q N1N438 VDD VDD pch W=6.3U L=0.24U
M10 Q N1N438 GVSS 0 nch W=3.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or4s3 Q DIN1 DIN2 DIN3 DIN4
M1 N1N425 DIN1 VDD VDD pch W=4.4U L=0.24U
M2 N1N441 DIN2 N1N425 VDD pch W=3.9U L=0.24U
M3 N1N441 DIN1 GVSS 0 nch W=1.7U L=0.24U
M4 N1N441 DIN2 GVSS 0 nch W=1.7U L=0.24U
M5 N1N422 DIN3 VDD VDD pch W=4.4U L=0.24U
M6 N1N428 DIN4 N1N422 VDD pch W=3.9U L=0.24U
M7 N1N428 DIN3 GVSS 0 nch W=1.7U L=0.24U
M8 N1N428 DIN4 GVSS 0 nch W=1.7U L=0.24U
M9 Q N1N441 VDD VDD pch W=4.2U L=0.24U
M11 Q N1N441 N1N445 0 nch W=4.2U L=0.24U
M12 N1N445 N1N428 GVSS 0 nch W=4.2U L=0.24U
M10 VDD N1N428 Q VDD pch W=4.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or5s1 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 GVSS 0 nch W=0.7U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=3U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=2.6U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=2.4U L=0.24U
M4 N1N444 DIN3 GVSS 0 nch W=0.7U L=0.24U
M6 N1N444 DIN1 GVSS 0 nch W=0.7U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=1.9U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=1.7U L=0.24U
M9 N1N494 DIN5 GVSS 0 nch W=0.7U L=0.24U
M10 GVSS DIN4 N1N494 0 nch W=0.7U L=0.24U
M11 Q N1N444 VDD VDD pch W=2U L=0.24U
M12 VDD N1N494 Q VDD pch W=2U L=0.24U
M13 Q N1N444 N1N480 0 nch W=1.7U L=0.24U
M14 N1N480 N1N494 GVSS 0 nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or5s2 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 GVSS 0 nch W=1.4U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=6U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=5.8U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=5.6U L=0.24U
M4 N1N444 DIN3 GVSS 0 nch W=1.4U L=0.24U
M6 N1N444 DIN1 GVSS 0 nch W=1.4U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=3.9U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=3.7U L=0.24U
M9 N1N494 DIN5 GVSS 0 nch W=1.4U L=0.24U
M10 GVSS DIN4 N1N494 0 nch W=1.4U L=0.24U
M11 Q N1N444 VDD VDD pch W=4U L=0.24U
M12 VDD N1N494 Q VDD pch W=4U L=0.24U
M13 Q N1N444 N1N480 0 nch W=3.6U L=0.24U
M14 N1N480 N1N494 GVSS 0 nch W=3.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_or5s3 Q DIN1 DIN2 DIN3 DIN4 DIN5
M5 N1N444 DIN2 GVSS 0 nch W=2.3U L=0.24U
M1 N1N440 DIN1 VDD VDD pch W=10.6U L=0.24U
M2 N1N442 DIN2 N1N440 VDD pch W=9.9U L=0.24U
M3 N1N444 DIN3 N1N442 VDD pch W=9.4U L=0.24U
M4 N1N444 DIN3 GVSS 0 nch W=2.3U L=0.24U
M6 N1N444 DIN1 GVSS 0 nch W=2.3U L=0.24U
M7 N1N489 DIN4 VDD VDD pch W=6.34U L=0.24U
M8 N1N494 DIN5 N1N489 VDD pch W=6.2U L=0.24U
M9 N1N494 DIN5 GVSS 0 nch W=2.3U L=0.24U
M10 GVSS DIN4 N1N494 0 nch W=2.3U L=0.24U
M11 Q N1N444 VDD VDD pch W=6.8U L=0.24U
M12 VDD N1N494 Q VDD pch W=6.8U L=0.24U
M13 Q N1N444 N1N480 0 nch W=5.7U L=0.24U
M14 N1N480 N1N494 GVSS 0 nch W=5.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ppt1s1 OUTD DIN OUTS
M1 OUTD DIN OUTS VDD pch W=2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ppt1s2 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ppt1s3 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ppt1s4 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ppt1s5 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=32U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ppt1s6 DIN OUTD OUTS
M1 OUTD DIN OUTS VDD pch W=64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ppu1s1 OUTD GIN
M1 OUTD GIN VDD VDD pch W=1.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ppu1s2 OUTD GIN
M1 OUTD GIN VDD VDD pch W=3.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_rpc1s1 DIN
M1 N1N254 N1N294 VDD VDD pch W=0.8U L=0.24U
M3 DIN N1N294 N1N258 0 nch W=0.8U L=0.24U
M2 DIN N1N294 N1N254 VDD pch W=0.8U L=0.24U
M4 N1N258 N1N294 GVSS 0 nch W=0.8U L=0.24U
M5 N1N294 DIN VDD VDD pch W=1.6U L=0.24U
M6 N1N294 DIN GVSS 0 nch W=1.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_rpc1s2 DIN
M1 N1N254 N1N294 VDD VDD pch W=1.2U L=0.24U
M3 DIN N1N294 N1N258 0 nch W=1.2U L=0.24U
M2 DIN N1N294 N1N254 VDD pch W=1.2U L=0.24U
M4 N1N258 N1N294 GVSS 0 nch W=1.2U L=0.24U
M5 N1N294 DIN VDD VDD pch W=2.5U L=0.24U
M6 N1N294 DIN GVSS 0 nch W=1.7U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffacs1 Q QN CLRB CLK SSEL SDIN DIN
M23 TP7 CLRB VDD VDD pch W=1.3U L=0.24U
M27 Q TP8 VDD VDD pch W=3.14U L=0.24U
M15 TP5 TP3 VDD VDD pch W=1.3U L=0.24U
M30 QN Q GVSS 0 nch W=1.42U L=0.24U
M9 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M10 TP21 TP1 TP3 0 nch W=0.8U L=0.24U
M19 TP5 CLK TP8 0 nch W=0.96U L=0.24U
M20 TP8 TP1 TP5 VDD pch W=1.4U L=0.24U
M12 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M21 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M22 TP8 TP1 TP7 0 nch W=0.8U L=0.24U
M29 QN Q VDD VDD pch W=3.02U L=0.24U
M11 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M17 TP5 TP3 TP6 0 nch W=0.9U L=0.24U
M25 TP7 Q TP9 0 nch W=0.9U L=0.24U
M28 Q TP8 GVSS 0 nch W=1.96U L=0.24U
M16 TP5 CLRB VDD VDD pch W=1.3U L=0.24U
M14 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M18 TP6 CLRB GVSS 0 nch W=0.9U L=0.24U
M7 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M24 TP7 Q VDD VDD pch W=1.3U L=0.24U
M26 TP9 CLRB GVSS 0 nch W=0.9U L=0.24U
M8 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffacs2 Q QN CLRB CLK SSEL SDIN DIN
M23 TP7 CLRB VDD VDD pch W=1.3U L=0.24U
M27 Q TP8 VDD VDD pch W=6.2U L=0.24U
M15 TP5 TP3 VDD VDD pch W=1.84U L=0.24U
M30 QN Q GVSS 0 nch W=2.68U L=0.24U
M9 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M10 TP21 TP1 TP3 0 nch W=0.8U L=0.24U
M19 TP5 CLK TP8 0 nch W=1.52U L=0.24U
M20 TP8 TP1 TP5 VDD pch W=1.9U L=0.24U
M12 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M21 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M22 TP8 TP1 TP7 0 nch W=0.8U L=0.24U
M29 QN Q VDD VDD pch W=6.16U L=0.24U
M11 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M17 TP5 TP3 TP6 0 nch W=1.48U L=0.24U
M25 TP7 Q TP9 0 nch W=0.9U L=0.24U
M28 Q TP8 GVSS 0 nch W=3.98U L=0.24U
M16 TP5 CLRB VDD VDD pch W=1.84U L=0.24U
M14 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M18 TP6 CLRB GVSS 0 nch W=1.48U L=0.24U
M7 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M13 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M24 TP7 Q VDD VDD pch W=1.3U L=0.24U
M26 TP9 CLRB GVSS 0 nch W=0.9U L=0.24U
M8 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffascs1 SETB CLRB DIN SSEL SDIN CLK QN Q
M18 TP6 CLK GVSS 0 nch W=0.8U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M12 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
M8 TP1 CLRB GVSS 0 nch W=0.8U L=0.24U
M7 TP1 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP1 VDD VDD pch W=2.2U L=0.24U
M10 TP4 TP1 GVSS 0 nch W=1.4U L=0.24U
M39 Q TP13 VDD VDD pch W=3.18U L=0.24U
M29 TP11 TP8 TP12 0 nch W=2.2U L=0.24U
M19 TP8 CLK TP21 VDD pch W=1.3U L=0.24U
M20 TP21 TP6 TP8 0 nch W=0.8U L=0.24U
M31 TP11 CLK TP13 0 nch W=2.2U L=0.24U
M32 TP13 TP6 TP11 VDD pch W=2.5U L=0.24U
M21 TP8 CLK TP9 0 nch W=0.8U L=0.24U
M22 TP9 TP6 TP8 VDD pch W=1.3U L=0.24U
M33 TP14 CLK TP13 VDD pch W=1.3U L=0.24U
M27 TP11 TP8 VDD VDD pch W=2.4U L=0.24U
M28 TP11 TP4 VDD VDD pch W=2.4U L=0.24U
M26 TP10 TP11 GVSS 0 nch W=0.8U L=0.24U
M38 TP15 TP4 GVSS 0 nch W=0.8U L=0.24U
M30 TP12 TP4 GVSS 0 nch W=2.2U L=0.24U
M42 TP16 TP13 GVSS 0 nch W=2.64U L=0.24U
M40 Q TP2 VDD VDD pch W=3.18U L=0.24U
M41 Q TP2 TP16 0 nch W=2.64U L=0.24U
M25 TP9 TP2 TP10 0 nch W=0.8U L=0.24U
M17 TP6 CLK VDD VDD pch W=1.4U L=0.24U
M15 TP2 TP0 TP3 0 nch W=1.3U L=0.24U
M16 TP3 TP4 GVSS 0 nch W=1.3U L=0.24U
M44 QN Q GVSS 0 nch W=1.44U L=0.24U
M13 TP2 TP0 VDD VDD pch W=1.8U L=0.24U
M14 TP2 TP4 VDD VDD pch W=1.8U L=0.24U
M23 TP9 TP2 VDD VDD pch W=1.3U L=0.24U
M24 TP9 TP11 VDD VDD pch W=1.3U L=0.24U
M37 TP14 Q TP15 0 nch W=0.8U L=0.24U
M36 TP14 Q VDD VDD pch W=1.3U L=0.24U
M34 TP13 TP6 TP14 0 nch W=0.8U L=0.24U
M43 QN Q VDD VDD pch W=3.18U L=0.24U
M11 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M35 TP14 TP4 VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffascs2 SETB CLRB DIN SSEL SDIN CLK QN Q
M18 TP6 CLK GVSS 0 nch W=0.8U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M12 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
M8 TP1 CLRB GVSS 0 nch W=0.8U L=0.24U
M7 TP1 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP4 TP1 VDD VDD pch W=2.7U L=0.24U
M10 TP4 TP1 GVSS 0 nch W=2.2U L=0.24U
M39 Q TP13 VDD VDD pch W=6.26U L=0.24U
M29 TP11 TP8 TP12 0 nch W=2.92U L=0.24U
M19 TP8 CLK TP21 VDD pch W=1.3U L=0.24U
M20 TP21 TP6 TP8 0 nch W=0.8U L=0.24U
M31 TP11 CLK TP13 0 nch W=2.7U L=0.24U
M32 TP13 TP6 TP11 VDD pch W=3U L=0.24U
M21 TP8 CLK TP9 0 nch W=0.8U L=0.24U
M22 TP9 TP6 TP8 VDD pch W=1.3U L=0.24U
M33 TP14 CLK TP13 VDD pch W=1.3U L=0.24U
M27 TP11 TP8 VDD VDD pch W=3.24U L=0.24U
M28 TP11 TP4 VDD VDD pch W=3.24U L=0.24U
M26 TP10 TP11 GVSS 0 nch W=0.8U L=0.24U
M38 TP15 TP4 GVSS 0 nch W=0.8U L=0.24U
M30 TP12 TP4 GVSS 0 nch W=2.92U L=0.24U
M42 TP16 TP13 GVSS 0 nch W=5.26U L=0.24U
M40 Q TP2 VDD VDD pch W=6.26U L=0.24U
M41 Q TP2 TP16 0 nch W=5.26U L=0.24U
M25 TP9 TP2 TP10 0 nch W=0.8U L=0.24U
M17 TP6 CLK VDD VDD pch W=1.6U L=0.24U
M15 TP2 TP0 TP3 0 nch W=2.2U L=0.24U
M16 TP3 TP4 GVSS 0 nch W=2.2U L=0.24U
M44 QN Q GVSS 0 nch W=2.88U L=0.24U
M13 TP2 TP0 VDD VDD pch W=2.82U L=0.24U
M14 TP2 TP4 VDD VDD pch W=2.82U L=0.24U
M23 TP9 TP2 VDD VDD pch W=1.3U L=0.24U
M24 TP9 TP11 VDD VDD pch W=1.3U L=0.24U
M37 TP14 Q TP15 0 nch W=0.8U L=0.24U
M36 TP14 Q VDD VDD pch W=1.3U L=0.24U
M34 TP13 TP6 TP14 0 nch W=0.8U L=0.24U
M43 QN Q VDD VDD pch W=6.2U L=0.24U
M11 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M35 TP14 TP4 VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffass1 Q QN SETB CLK SSEL SDIN DIN
M27 TP7 SETB VDD VDD pch W=1.3U L=0.24U
M19 TP5 TP3 VDD VDD pch W=1.3U L=0.24U
M34 Q QN GVSS 0 nch W=1.42U L=0.24U
M13 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M14 TP21 TP1 TP3 0 nch W=0.8U L=0.24U
M23 TP5 CLK TP8 0 nch W=0.96U L=0.24U
M24 TP8 TP1 TP5 VDD pch W=1.4U L=0.24U
M16 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M25 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M33 Q QN VDD VDD pch W=3.02U L=0.24U
M15 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M29 TP7 QN TP9 0 nch W=0.9U L=0.24U
M32 QN TP8 GVSS 0 nch W=1.96U L=0.24U
M20 TP5 SETB VDD VDD pch W=1.3U L=0.24U
M18 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M22 TP6 SETB GVSS 0 nch W=0.9U L=0.24U
M17 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M30 TP9 SETB GVSS 0 nch W=0.9U L=0.24U
M28 TP7 QN VDD VDD pch W=1.3U L=0.24U
M21 TP5 TP3 TP6 0 nch W=0.9U L=0.24U
M12 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M26 TP8 TP1 TP7 0 nch W=0.8U L=0.24U
M31 QN TP8 VDD VDD pch W=3.14U L=0.24U
M11 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M3 TP19 SDIN VDD VDD pch W=1.3U L=0.24U
M4 TP19 SDIN GVSS 0 nch W=0.8U L=0.24U
M1 TP18 DIN VDD VDD pch W=1.3U L=0.24U
M2 TP18 DIN GVSS 0 nch W=0.8U L=0.24U
M9 TP21 TP20 TP19 VDD pch W=1.3U L=0.24U
M10 TP19 SSEL TP21 0 nch W=0.8U L=0.24U
M5 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M6 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M8 TP18 TP20 TP21 0 nch W=0.8U L=0.24U
M7 TP21 SSEL TP18 VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffass2 Q QN SETB CLK SSEL SDIN DIN
M27 TP7 SETB VDD VDD pch W=1.3U L=0.24U
M19 TP5 TP3 VDD VDD pch W=1.84U L=0.24U
M34 Q QN GVSS 0 nch W=2.68U L=0.24U
M13 TP3 CLK TP21 VDD pch W=1.3U L=0.24U
M14 TP21 TP1 TP3 0 nch W=0.8U L=0.24U
M23 TP5 CLK TP8 0 nch W=1.52U L=0.24U
M24 TP8 TP1 TP5 VDD pch W=1.9U L=0.24U
M16 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M25 TP7 CLK TP8 VDD pch W=1.3U L=0.24U
M33 Q QN VDD VDD pch W=6.16U L=0.24U
M15 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M29 TP7 QN TP9 0 nch W=0.9U L=0.24U
M32 QN TP8 GVSS 0 nch W=3.98U L=0.24U
M20 TP5 SETB VDD VDD pch W=1.84U L=0.24U
M18 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M22 TP6 SETB GVSS 0 nch W=1.48U L=0.24U
M17 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M30 TP9 SETB GVSS 0 nch W=0.9U L=0.24U
M28 TP7 QN VDD VDD pch W=1.3U L=0.24U
M21 TP5 TP3 TP6 0 nch W=1.48U L=0.24U
M12 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M26 TP8 TP1 TP7 0 nch W=0.8U L=0.24U
M31 QN TP8 VDD VDD pch W=6.2U L=0.24U
M11 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M3 TP19 SDIN VDD VDD pch W=1.3U L=0.24U
M4 TP19 SDIN GVSS 0 nch W=0.8U L=0.24U
M1 TP18 DIN VDD VDD pch W=1.3U L=0.24U
M2 TP18 DIN GVSS 0 nch W=0.8U L=0.24U
M9 TP21 TP20 TP19 VDD pch W=1.3U L=0.24U
M10 TP19 SSEL TP21 0 nch W=0.8U L=0.24U
M5 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M6 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M8 TP18 TP20 TP21 0 nch W=0.8U L=0.24U
M7 TP21 SSEL TP18 VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffcs1 SSEL CLRB DIN SDIN CLK Q QN
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M9 TP2 TP21 TP1 0 nch W=0.8U L=0.24U
M8 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M7 TP2 TP21 VDD VDD pch W=1.3U L=0.24U
M12 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M13 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M14 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M19 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M21 TP6 CLK TP7 0 nch W=0.8U L=0.24U
M22 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M27 QN TP7 VDD VDD pch W=3.14U L=0.24U
M28 QN TP7 GVSS 0 nch W=2.06U L=0.24U
M15 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M16 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M18 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M23 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M29 Q QN VDD VDD pch W=2.94U L=0.24U
M30 Q QN GVSS 0 nch W=1.28U L=0.24U
M20 TP6 TP4 GVSS 0 nch W=0.8U L=0.24U
M11 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M26 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M24 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M25 TP8 QN VDD VDD pch W=1.3U L=0.24U
M17 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M10 TP1 CLRB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffcs2 SSEL CLRB DIN SDIN CLK Q QN
M13 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M14 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M19 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M21 TP6 CLK TP7 0 nch W=1.3U L=0.24U
M22 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M27 QN TP7 VDD VDD pch W=6.24U L=0.24U
M28 QN TP7 GVSS 0 nch W=3.98U L=0.24U
M15 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M16 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M17 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M18 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M23 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M24 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M25 TP8 QN VDD VDD pch W=1.3U L=0.24U
M26 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M29 Q QN VDD VDD pch W=5.92U L=0.24U
M30 Q QN GVSS 0 nch W=2.66U L=0.24U
M20 TP6 TP4 GVSS 0 nch W=1.26U L=0.24U
M11 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M12 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M7 TP2 TP21 VDD VDD pch W=1.3U L=0.24U
M8 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M9 TP2 TP21 TP1 0 nch W=0.8U L=0.24U
M10 TP1 CLRB GVSS 0 nch W=0.8U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffles1 EB DIN SSEL SDIN CLK QN Q
M29 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M30 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M40 TP9 TP10 GVSS 0 nch W=0.8U L=0.24U
M50 Q TP11 GVSS 0 nch W=2.06U L=0.24U
M42 TP10 TP8 GVSS 0 nch W=0.8U L=0.24U
M48 TP5 Q GVSS 0 nch W=0.8U L=0.24U
M47 TP5 Q VDD VDD pch W=1.3U L=0.24U
M52 QN Q GVSS 0 nch W=1.28U L=0.24U
M35 TP8 CLK TP3 VDD pch W=1.3U L=0.24U
M36 TP3 TP7 TP8 0 nch W=0.8U L=0.24U
M43 TP10 CLK TP11 0 nch W=0.8U L=0.24U
M38 TP9 TP7 TP8 VDD pch W=1.3U L=0.24U
M46 TP11 TP7 TP5 0 nch W=0.8U L=0.24U
M51 QN Q VDD VDD pch W=2.94U L=0.24U
M37 TP8 CLK TP9 0 nch W=0.8U L=0.24U
M49 Q TP11 VDD VDD pch W=3.14U L=0.24U
M41 TP10 TP8 VDD VDD pch W=1.8U L=0.24U
M39 TP9 TP10 VDD VDD pch W=1.3U L=0.24U
M44 TP11 TP7 TP10 VDD pch W=1.3U L=0.24U
M45 TP5 CLK TP11 VDD pch W=1.3U L=0.24U
M19 TP3 TP23 SDIN VDD pch W=1.3U L=0.24U
M20 SDIN SSEL TP3 0 nch W=0.8U L=0.24U
M28 TP27 TP25 GVSS 0 nch W=0.8U L=0.24U
M27 TP27 TP25 VDD VDD pch W=1.3U L=0.24U
M21 TP25 EB VDD VDD pch W=1.3U L=0.24U
M23 TP25 EB TP26 0 nch W=0.8U L=0.24U
M24 TP26 TP23 GVSS 0 nch W=0.8U L=0.24U
M6 TP22 TP23 GVSS 0 nch W=0.8U L=0.24U
M18 TP24 TP21 GVSS 0 nch W=0.8U L=0.24U
M17 TP24 TP21 VDD VDD pch W=1.3U L=0.24U
M3 TP21 TP20 VDD VDD pch W=1.3U L=0.24U
M5 TP21 TP20 TP22 0 nch W=0.8U L=0.24U
M2 TP20 EB GVSS 0 nch W=0.8U L=0.24U
M1 TP20 EB VDD VDD pch W=1.3U L=0.24U
M15 TP3 TP21 DIN VDD pch W=1.3U L=0.24U
M16 DIN TP24 TP3 0 nch W=0.8U L=0.24U
M25 TP4 TP25 TP3 VDD pch W=1.3U L=0.24U
M26 TP3 TP27 TP4 0 nch W=0.8U L=0.24U
M4 TP21 TP23 VDD VDD pch W=1.3U L=0.24U
M22 TP25 TP23 VDD VDD pch W=1.3U L=0.24U
M34 TP7 CLK GVSS 0 nch W=0.8U L=0.24U
M33 TP7 CLK VDD VDD pch W=1.3U L=0.24U
M11 TP23 SSEL VDD VDD pch W=1.5U L=0.24U
M12 TP23 SSEL GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffles2 EB DIN SSEL SDIN CLK QN Q
M29 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M30 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M40 TP9 TP10 GVSS 0 nch W=0.8U L=0.24U
M50 Q TP11 GVSS 0 nch W=3.98U L=0.24U
M42 TP10 TP8 GVSS 0 nch W=1.26U L=0.24U
M48 TP5 Q GVSS 0 nch W=0.8U L=0.24U
M47 TP5 Q VDD VDD pch W=1.3U L=0.24U
M52 QN Q GVSS 0 nch W=2.66U L=0.24U
M35 TP8 CLK TP3 VDD pch W=1.3U L=0.24U
M36 TP3 TP7 TP8 0 nch W=0.8U L=0.24U
M43 TP10 CLK TP11 0 nch W=1.3U L=0.24U
M38 TP9 TP7 TP8 VDD pch W=1.3U L=0.24U
M46 TP11 TP7 TP5 0 nch W=0.8U L=0.24U
M51 QN Q VDD VDD pch W=5.92U L=0.24U
M37 TP8 CLK TP9 0 nch W=0.8U L=0.24U
M49 Q TP11 VDD VDD pch W=6.24U L=0.24U
M41 TP10 TP8 VDD VDD pch W=2.78U L=0.24U
M39 TP9 TP10 VDD VDD pch W=1.3U L=0.24U
M44 TP11 TP7 TP10 VDD pch W=1.8U L=0.24U
M45 TP5 CLK TP11 VDD pch W=1.3U L=0.24U
M19 TP3 TP23 SDIN VDD pch W=1.3U L=0.24U
M20 SDIN SSEL TP3 0 nch W=0.8U L=0.24U
M28 TP27 TP25 GVSS 0 nch W=0.8U L=0.24U
M27 TP27 TP25 VDD VDD pch W=1.3U L=0.24U
M21 TP25 EB VDD VDD pch W=1.3U L=0.24U
M23 TP25 EB TP26 0 nch W=0.8U L=0.24U
M24 TP26 TP23 GVSS 0 nch W=0.8U L=0.24U
M6 TP22 TP23 GVSS 0 nch W=0.8U L=0.24U
M18 TP24 TP21 GVSS 0 nch W=0.8U L=0.24U
M17 TP24 TP21 VDD VDD pch W=1.3U L=0.24U
M3 TP21 TP20 VDD VDD pch W=1.3U L=0.24U
M5 TP21 TP20 TP22 0 nch W=0.8U L=0.24U
M2 TP20 EB GVSS 0 nch W=0.8U L=0.24U
M1 TP20 EB VDD VDD pch W=1.3U L=0.24U
M15 TP3 TP21 DIN VDD pch W=1.3U L=0.24U
M16 DIN TP24 TP3 0 nch W=0.8U L=0.24U
M25 TP4 TP25 TP3 VDD pch W=1.3U L=0.24U
M26 TP3 TP27 TP4 0 nch W=0.8U L=0.24U
M4 TP21 TP23 VDD VDD pch W=1.3U L=0.24U
M22 TP25 TP23 VDD VDD pch W=1.3U L=0.24U
M34 TP7 CLK GVSS 0 nch W=0.8U L=0.24U
M33 TP7 CLK VDD VDD pch W=1.3U L=0.24U
M11 TP23 SSEL VDD VDD pch W=1.5U L=0.24U
M12 TP23 SSEL GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffs1 Q QN CLK SSEL SDIN DIN
M17 TP3 CLK TP9 VDD pch W=1.3U L=0.24U
M18 TP9 TP1 TP3 0 nch W=0.8U L=0.24U
M21 TP5 TP3 VDD VDD pch W=1.8U L=0.24U
M25 TP5 CLK TP6 0 nch W=0.8U L=0.24U
M26 TP6 TP1 TP5 VDD pch W=1.3U L=0.24U
M29 Q TP6 VDD VDD pch W=3.14U L=0.24U
M30 Q TP6 GVSS 0 nch W=2.06U L=0.24U
M19 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M20 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M23 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M24 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M27 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M28 TP6 TP1 TP7 0 nch W=0.8U L=0.24U
M31 TP7 Q VDD VDD pch W=1.3U L=0.24U
M32 TP7 Q GVSS 0 nch W=0.8U L=0.24U
M33 QN Q VDD VDD pch W=2.94U L=0.24U
M34 QN Q GVSS 0 nch W=1.28U L=0.24U
M22 TP5 TP3 GVSS 0 nch W=0.8U L=0.24U
M14 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M13 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M9 DIN TP8 TP9 0 nch W=0.8U L=0.24U
M10 TP9 SSEL DIN VDD pch W=1.3U L=0.24U
M11 TP9 TP8 SDIN VDD pch W=1.3U L=0.24U
M12 SDIN SSEL TP9 0 nch W=0.8U L=0.24U
M6 TP8 SSEL GVSS 0 nch W=0.8U L=0.24U
M5 TP8 SSEL VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffs2 Q QN CLK SSEL SDIN DIN
M17 TP3 CLK TP9 VDD pch W=1.3U L=0.24U
M18 TP9 TP1 TP3 0 nch W=0.8U L=0.24U
M21 TP5 TP3 VDD VDD pch W=2.76U L=0.24U
M25 TP5 CLK TP6 0 nch W=1.3U L=0.24U
M26 TP6 TP1 TP5 VDD pch W=1.8U L=0.24U
M29 Q TP6 VDD VDD pch W=6.24U L=0.24U
M30 Q TP6 GVSS 0 nch W=3.98U L=0.24U
M19 TP3 CLK TP4 0 nch W=0.8U L=0.24U
M20 TP4 TP1 TP3 VDD pch W=1.3U L=0.24U
M23 TP4 TP5 VDD VDD pch W=1.3U L=0.24U
M24 TP4 TP5 GVSS 0 nch W=0.8U L=0.24U
M27 TP7 CLK TP6 VDD pch W=1.3U L=0.24U
M28 TP6 TP1 TP7 0 nch W=0.8U L=0.24U
M31 TP7 Q VDD VDD pch W=1.3U L=0.24U
M32 TP7 Q GVSS 0 nch W=0.8U L=0.24U
M33 QN Q VDD VDD pch W=5.92U L=0.24U
M34 QN Q GVSS 0 nch W=2.66U L=0.24U
M22 TP5 TP3 GVSS 0 nch W=1.26U L=0.24U
M14 TP1 CLK GVSS 0 nch W=0.8U L=0.24U
M13 TP1 CLK VDD VDD pch W=1.3U L=0.24U
M9 DIN TP8 TP9 0 nch W=0.8U L=0.24U
M10 TP9 SSEL DIN VDD pch W=1.3U L=0.24U
M11 TP9 TP8 SDIN VDD pch W=1.3U L=0.24U
M12 SDIN SSEL TP9 0 nch W=0.8U L=0.24U
M6 TP8 SSEL GVSS 0 nch W=0.8U L=0.24U
M5 TP8 SSEL VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffscs1 SSEL CLR DIN SET SDIN CLK QN Q
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M17 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M18 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M23 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M25 TP6 CLK TP7 0 nch W=0.8U L=0.24U
M26 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M31 QN TP7 VDD VDD pch W=3.14U L=0.24U
M32 QN TP7 GVSS 0 nch W=2.06U L=0.24U
M19 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M20 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M22 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M27 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M33 Q QN VDD VDD pch W=2.94U L=0.24U
M34 Q QN GVSS 0 nch W=1.28U L=0.24U
M24 TP6 TP4 GVSS 0 nch W=0.8U L=0.24U
M15 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M16 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M30 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M28 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M29 TP8 QN VDD VDD pch W=1.3U L=0.24U
M21 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M9 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M10 TP2 TP21 TP1 VDD pch W=1.3U L=0.24U
M11 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M12 TP2 CLRB TP9 0 nch W=0.8U L=0.24U
M13 TP9 TP21 GVSS 0 nch W=0.8U L=0.24U
M14 TP9 TP0 GVSS 0 nch W=0.8U L=0.24U
M7 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M8 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffscs2 SSEL CLR DIN SET SDIN CLK QN Q
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M17 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M18 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M23 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M25 TP6 CLK TP7 0 nch W=1.3U L=0.24U
M26 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M31 QN TP7 VDD VDD pch W=6.24U L=0.24U
M32 QN TP7 GVSS 0 nch W=3.98U L=0.24U
M19 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M20 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M22 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M27 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M33 Q QN VDD VDD pch W=5.92U L=0.24U
M34 Q QN GVSS 0 nch W=2.66U L=0.24U
M24 TP6 TP4 GVSS 0 nch W=1.26U L=0.24U
M15 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M16 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M30 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M28 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M29 TP8 QN VDD VDD pch W=1.3U L=0.24U
M21 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M9 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M10 TP2 TP21 TP1 VDD pch W=1.3U L=0.24U
M11 TP2 CLRB VDD VDD pch W=1.3U L=0.24U
M12 TP2 CLRB TP9 0 nch W=0.8U L=0.24U
M13 TP9 TP21 GVSS 0 nch W=0.8U L=0.24U
M14 TP9 TP0 GVSS 0 nch W=0.8U L=0.24U
M7 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M8 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffss1 SETB DIN SSEL SDIN CLK QN Q
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M8 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
M7 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M14 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M15 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M16 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M21 TP6 TP4 VDD VDD pch W=1.8U L=0.24U
M23 TP6 CLK TP7 0 nch W=0.8U L=0.24U
M24 TP7 TP3 TP6 VDD pch W=1.3U L=0.24U
M29 QN TP7 VDD VDD pch W=3.14U L=0.24U
M30 QN TP7 GVSS 0 nch W=2.06U L=0.24U
M17 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M18 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M20 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M25 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M31 Q QN VDD VDD pch W=2.94U L=0.24U
M32 Q QN GVSS 0 nch W=1.28U L=0.24U
M22 TP6 TP4 GVSS 0 nch W=0.8U L=0.24U
M13 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M28 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M11 TP2 TP21 GVSS 0 nch W=0.8U L=0.24U
M12 TP2 TP0 GVSS 0 nch W=0.8U L=0.24U
M26 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M27 TP8 QN VDD VDD pch W=1.3U L=0.24U
M19 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M9 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M10 TP2 TP21 TP1 VDD pch W=1.3U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sdffss2 SETB DIN SSEL SDIN CLK QN Q
M6 SDIN SSEL TP21 0 nch W=0.8U L=0.24U
M3 TP21 SSEL DIN VDD pch W=1.3U L=0.24U
M8 TP0 SETB GVSS 0 nch W=0.8U L=0.24U
M7 TP0 SETB VDD VDD pch W=1.3U L=0.24U
M14 TP3 CLK GVSS 0 nch W=0.8U L=0.24U
M15 TP4 CLK TP2 VDD pch W=1.3U L=0.24U
M16 TP2 TP3 TP4 0 nch W=0.8U L=0.24U
M21 TP6 TP4 VDD VDD pch W=2.76U L=0.24U
M23 TP6 CLK TP7 0 nch W=1.3U L=0.24U
M24 TP7 TP3 TP6 VDD pch W=1.8U L=0.24U
M29 QN TP7 VDD VDD pch W=6.24U L=0.24U
M30 QN TP7 GVSS 0 nch W=3.98U L=0.24U
M17 TP4 CLK TP5 0 nch W=0.8U L=0.24U
M18 TP5 TP3 TP4 VDD pch W=1.3U L=0.24U
M20 TP5 TP6 GVSS 0 nch W=0.8U L=0.24U
M25 TP8 CLK TP7 VDD pch W=1.3U L=0.24U
M31 Q QN VDD VDD pch W=5.92U L=0.24U
M32 Q QN GVSS 0 nch W=2.66U L=0.24U
M22 TP6 TP4 GVSS 0 nch W=1.26U L=0.24U
M13 TP3 CLK VDD VDD pch W=1.3U L=0.24U
M28 TP8 QN GVSS 0 nch W=0.8U L=0.24U
M11 TP2 TP21 GVSS 0 nch W=0.8U L=0.24U
M12 TP2 TP0 GVSS 0 nch W=0.8U L=0.24U
M26 TP7 TP3 TP8 0 nch W=0.8U L=0.24U
M27 TP8 QN VDD VDD pch W=1.3U L=0.24U
M19 TP5 TP6 VDD VDD pch W=1.3U L=0.24U
M1 TP20 SSEL VDD VDD pch W=1.3U L=0.24U
M2 TP20 SSEL GVSS 0 nch W=0.8U L=0.24U
M4 DIN TP20 TP21 0 nch W=0.8U L=0.24U
M9 TP1 TP0 VDD VDD pch W=1.3U L=0.24U
M10 TP2 TP21 TP1 VDD pch W=1.3U L=0.24U
M5 TP21 TP20 SDIN VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sub1s1 OUTD OUTC0 AIN BIN CIN
M5 N1N303 N1N388 N1N305 0 nch W=0.8U L=0.24U
M3 N1N301 AIN VDD VDD pch W=1.2U L=0.24U
M4 N1N303 N1N388 N1N301 VDD pch W=1.1U L=0.24U
M7 N1N307 AIN VDD VDD pch W=1.2U L=0.24U
M8 VDD N1N388 N1N307 VDD pch W=1.2U L=0.24U
M9 N1N307 CIN N1N303 VDD pch W=1.1U L=0.24U
M6 N1N305 AIN GVSS 0 nch W=0.9U L=0.24U
M10 N1N312 CIN N1N303 0 nch W=0.8U L=0.24U
M12 GVSS N1N388 N1N312 0 nch W=0.9U L=0.24U
M11 N1N312 AIN GVSS 0 nch W=0.9U L=0.24U
M13 N1N337 AIN VDD VDD pch W=1.4U L=0.24U
M17 N1N341 N1N303 N1N337 VDD pch W=1.1U L=0.24U
M14 VDD CIN N1N337 VDD pch W=1.4U L=0.24U
M18 N1N341 N1N303 N1N366 0 nch W=0.9U L=0.24U
M20 N1N366 CIN GVSS 0 nch W=0.9U L=0.24U
M19 N1N366 AIN GVSS 0 nch W=0.9U L=0.24U
M21 GVSS N1N388 N1N366 0 nch W=0.9U L=0.24U
M15 VDD N1N388 N1N337 VDD pch W=1.4U L=0.24U
M16 VDD AIN N1N359 VDD pch W=2.1U L=0.24U
M22 N1N359 N1N388 N1N357 VDD pch W=2.1U L=0.24U
M23 N1N357 CIN N1N341 VDD pch W=2.1U L=0.24U
M24 N1N348 CIN N1N341 0 nch W=1.3U L=0.24U
M25 N1N352 N1N388 N1N348 0 nch W=1.3U L=0.24U
M26 GVSS AIN N1N352 0 nch W=1.3U L=0.24U
M28 OUTD N1N341 GVSS 0 nch W=0.9U L=0.24U
M27 OUTD N1N341 VDD VDD pch W=1.36U L=0.24U
M2 N1N388 BIN GVSS 0 nch W=0.6U L=0.24U
M1 N1N388 BIN VDD VDD pch W=1.2U L=0.24U
M30 OUTC0 N1N303 GVSS 0 nch W=0.9U L=0.24U
M29 OUTC0 N1N303 VDD VDD pch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sub1s2 OUTD OUTC0 AIN BIN CIN
M5 N1N303 N1N388 N1N305 0 nch W=1.1U L=0.24U
M3 N1N301 AIN VDD VDD pch W=1.8U L=0.24U
M4 N1N303 N1N388 N1N301 VDD pch W=1.7U L=0.24U
M7 N1N307 AIN VDD VDD pch W=1.8U L=0.24U
M8 VDD N1N388 N1N307 VDD pch W=1.8U L=0.24U
M9 N1N307 CIN N1N303 VDD pch W=1.7U L=0.24U
M6 N1N305 AIN GVSS 0 nch W=1.2U L=0.24U
M10 N1N312 CIN N1N303 0 nch W=1.1U L=0.24U
M12 GVSS N1N388 N1N312 0 nch W=1.2U L=0.24U
M11 N1N312 AIN GVSS 0 nch W=1.2U L=0.24U
M13 N1N337 AIN VDD VDD pch W=2.1U L=0.24U
M17 N1N341 N1N303 N1N337 VDD pch W=1.66U L=0.24U
M14 VDD CIN N1N337 VDD pch W=2.1U L=0.24U
M18 N1N341 N1N303 N1N366 0 nch W=1.16U L=0.24U
M20 N1N366 CIN GVSS 0 nch W=1.16U L=0.24U
M19 N1N366 AIN GVSS 0 nch W=1.16U L=0.24U
M21 GVSS N1N388 N1N366 0 nch W=1.16U L=0.24U
M15 VDD N1N388 N1N337 VDD pch W=2.1U L=0.24U
M16 VDD AIN N1N359 VDD pch W=3.16U L=0.24U
M22 N1N359 N1N388 N1N357 VDD pch W=3.16U L=0.24U
M23 N1N357 CIN N1N341 VDD pch W=3.16U L=0.24U
M24 N1N348 CIN N1N341 0 nch W=1.74U L=0.24U
M25 N1N352 N1N388 N1N348 0 nch W=1.74U L=0.24U
M26 GVSS AIN N1N352 0 nch W=1.74U L=0.24U
M28 OUTD N1N341 GVSS 0 nch W=1.44U L=0.24U
M27 OUTD N1N341 VDD VDD pch W=2.48U L=0.24U
M2 N1N388 BIN GVSS 0 nch W=0.6U L=0.24U
M1 N1N388 BIN VDD VDD pch W=1.2U L=0.24U
M30 OUTC0 N1N303 GVSS 0 nch W=1.46U L=0.24U
M29 OUTC0 N1N303 VDD VDD pch W=2.32U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_sub1s3 OUTD OUTC0 AIN BIN CIN
M5 N1N303 N1N388 N1N305 0 nch W=1.6U L=0.24U
M3 N1N301 AIN VDD VDD pch W=2.7U L=0.24U
M4 N1N303 N1N388 N1N301 VDD pch W=2.6U L=0.24U
M7 N1N307 AIN VDD VDD pch W=2.7U L=0.24U
M8 VDD N1N388 N1N307 VDD pch W=2.7U L=0.24U
M9 N1N307 CIN N1N303 VDD pch W=2.6U L=0.24U
M6 N1N305 AIN GVSS 0 nch W=1.7U L=0.24U
M10 N1N312 CIN N1N303 0 nch W=1.6U L=0.24U
M12 GVSS N1N388 N1N312 0 nch W=1.7U L=0.24U
M11 N1N312 AIN GVSS 0 nch W=1.7U L=0.24U
M13 N1N337 AIN VDD VDD pch W=2.9U L=0.24U
M17 N1N341 N1N303 N1N337 VDD pch W=2.8U L=0.24U
M14 VDD CIN N1N337 VDD pch W=2.9U L=0.24U
M18 N1N341 N1N303 N1N366 0 nch W=1.52U L=0.24U
M20 N1N366 CIN GVSS 0 nch W=1.52U L=0.24U
M19 N1N366 AIN GVSS 0 nch W=1.52U L=0.24U
M21 GVSS N1N388 N1N366 0 nch W=1.52U L=0.24U
M15 VDD N1N388 N1N337 VDD pch W=2.9U L=0.24U
M16 VDD AIN N1N359 VDD pch W=4.4U L=0.24U
M22 N1N359 N1N388 N1N357 VDD pch W=4.4U L=0.24U
M23 N1N357 CIN N1N341 VDD pch W=4.3U L=0.24U
M24 N1N348 CIN N1N341 0 nch W=2.26U L=0.24U
M25 N1N352 N1N388 N1N348 0 nch W=2.26U L=0.24U
M26 GVSS AIN N1N352 0 nch W=2.26U L=0.24U
M28 OUTD N1N341 GVSS 0 nch W=2.9U L=0.24U
M27 OUTD N1N341 VDD VDD pch W=5U L=0.24U
M2 N1N388 BIN GVSS 0 nch W=0.7U L=0.24U
M1 N1N388 BIN VDD VDD pch W=1.4U L=0.24U
M30 OUTC0 N1N303 GVSS 0 nch W=2.9U L=0.24U
M29 OUTC0 N1N303 VDD VDD pch W=4.64U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibh1s1 Q E DIN
M2 N1N502 E GVSS 0 nch W=0.8U L=0.24U
M1 N1N502 E VDD VDD pch W=1.2U L=0.24U
M5 Q E N1N508 0 nch W=0.8U L=0.24U
M3 N1N504 DIN VDD VDD pch W=2.3U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=2.3U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibh1s2 Q E DIN
M2 N1N502 E GVSS 0 nch W=0.9U L=0.24U
M1 N1N502 E VDD VDD pch W=1.6U L=0.24U
M5 Q E N1N508 0 nch W=1U L=0.24U
M3 N1N504 DIN VDD VDD pch W=3U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=3U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibh1s3 Q E DIN
M2 N1N502 E GVSS 0 nch W=1.1U L=0.24U
M1 N1N502 E VDD VDD pch W=2.1U L=0.24U
M5 Q E N1N508 0 nch W=1.3U L=0.24U
M3 N1N504 DIN VDD VDD pch W=3.9U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=3.9U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibh1s4 Q E DIN
M2 N1N502 E GVSS 0 nch W=2U L=0.24U
M1 N1N502 E VDD VDD pch W=3U L=0.24U
M5 Q E N1N508 0 nch W=2.1U L=0.24U
M3 N1N504 DIN VDD VDD pch W=6.3U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=6.3U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=2.1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibh1s5 Q E DIN
M2 N1N502 E GVSS 0 nch W=2.3U L=0.24U
M1 N1N502 E VDD VDD pch W=3.7U L=0.24U
M5 Q E N1N508 0 nch W=3U L=0.24U
M3 N1N504 DIN VDD VDD pch W=9.32U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=9.32U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibh1s6 Q E DIN
M2 N1N502 E GVSS 0 nch W=2.9U L=0.24U
M1 N1N502 E VDD VDD pch W=4.8U L=0.24U
M3 N1N504 DIN VDD VDD pch W=11.4U L=0.24U
M4 Q N1N502 N1N504 VDD pch W=11.4U L=0.24U
M5 Q E N1N508 0 nch W=3.6U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=3.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibl1s1 Q EB DIN
M2 N1N510 EB GVSS 0 nch W=0.8U L=0.24U
M1 N1N510 EB VDD VDD pch W=1.2U L=0.24U
M3 N1N504 DIN VDD VDD pch W=2.2U L=0.24U
M4 Q EB N1N504 VDD pch W=2.2U L=0.24U
M5 Q N1N510 N1N508 0 nch W=0.86U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=0.86U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibl1s2 Q EB DIN
M2 N1N510 EB GVSS 0 nch W=0.9U L=0.24U
M1 N1N510 EB VDD VDD pch W=1.6U L=0.24U
M3 N1N504 DIN VDD VDD pch W=2.8U L=0.24U
M4 Q EB N1N504 VDD pch W=2.8U L=0.24U
M5 Q N1N510 N1N508 0 nch W=1.16U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=1.16U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibl1s3 Q EB DIN
M2 N1N510 EB GVSS 0 nch W=1.1U L=0.24U
M1 N1N510 EB VDD VDD pch W=2.1U L=0.24U
M3 N1N504 DIN VDD VDD pch W=3.6U L=0.24U
M4 Q EB N1N504 VDD pch W=3.6U L=0.24U
M5 Q N1N510 N1N508 0 nch W=1.5U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=1.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibl1s4 Q EB DIN
M2 N1N510 EB GVSS 0 nch W=1.8U L=0.24U
M1 N1N510 EB VDD VDD pch W=3.5U L=0.24U
M3 N1N504 DIN VDD VDD pch W=5.4U L=0.24U
M4 Q EB N1N504 VDD pch W=5.4U L=0.24U
M5 Q N1N510 N1N508 0 nch W=2.4U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=2.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibl1s5 Q EB DIN
M2 N1N510 EB GVSS 0 nch W=1.8U L=0.24U
M1 N1N510 EB VDD VDD pch W=3.7U L=0.24U
M3 N1N504 DIN VDD VDD pch W=8.7U L=0.24U
M4 Q EB N1N504 VDD pch W=8.7U L=0.24U
M5 Q N1N510 N1N508 0 nch W=4.5U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=4.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tibl1s6 Q EB DIN
M2 N1N510 EB GVSS 0 nch W=2.2U L=0.24U
M1 N1N510 EB VDD VDD pch W=4.4U L=0.24U
M3 N1N504 DIN VDD VDD pch W=11.3U L=0.24U
M4 Q EB N1N504 VDD pch W=11.3U L=0.24U
M5 Q N1N510 N1N508 0 nch W=6.2U L=0.24U
M6 N1N508 DIN GVSS 0 nch W=6.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbh1s1 Q E DIN
M2 N1N517 N1N509 VDD VDD pch W=2.6U L=0.24U
M1 N1N513 E VDD VDD pch W=1.5U L=0.24U
M4 N1N513 E GVSS 0 nch W=0.9U L=0.24U
M6 Q E N1N523 0 nch W=0.94U L=0.24U
M8 N1N523 N1N509 GVSS 0 nch W=0.94U L=0.24U
M7 N1N509 DIN GVSS 0 nch W=0.8U L=0.24U
M3 Q N1N513 N1N517 VDD pch W=2.6U L=0.24U
M5 N1N509 DIN VDD VDD pch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbh1s2 Q E DIN
M2 N1N286 E GVSS 0 nch W=0.9U L=0.24U
M1 N1N286 E VDD VDD pch W=1.6U L=0.24U
M4 N1N260 DIN GVSS 0 nch W=0.8U L=0.24U
M3 N1N260 DIN VDD VDD pch W=1.6U L=0.24U
M8 N1N267 N1N260 GVSS 0 nch W=1.24U L=0.24U
M7 Q E N1N267 0 nch W=1.24U L=0.24U
M6 Q N1N286 N1N262 VDD pch W=3.6U L=0.24U
M5 N1N262 N1N260 VDD VDD pch W=3.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbh1s3 Q E DIN
M6 N1N565 DIN VDD VDD pch W=1.4U L=0.24U
M1 N1N563 E VDD VDD pch W=1.3U L=0.24U
M3 N1N565 E VDD VDD pch W=1.4U L=0.24U
M9 Q N1N565 VDD VDD pch W=2.42U L=0.24U
M7 N1N567 N1N563 N1N565 VDD pch W=1.3U L=0.24U
M8 N1N567 DIN GVSS 0 nch W=0.9U L=0.24U
M10 Q N1N567 GVSS 0 nch W=1.46U L=0.24U
M4 N1N565 E N1N567 0 nch W=0.8U L=0.24U
M2 N1N563 E GVSS 0 nch W=0.8U L=0.24U
M5 N1N567 N1N563 GVSS 0 nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbh1s4 Q E DIN
M6 N1N565 DIN VDD VDD pch W=2.4U L=0.24U
M1 N1N563 E VDD VDD pch W=1.3U L=0.24U
M3 N1N565 E VDD VDD pch W=2U L=0.24U
M9 Q N1N565 VDD VDD pch W=3.3U L=0.24U
M7 N1N567 N1N563 N1N565 VDD pch W=2.6U L=0.24U
M8 N1N567 DIN GVSS 0 nch W=1.2U L=0.24U
M10 Q N1N567 GVSS 0 nch W=1.9U L=0.24U
M4 N1N565 E N1N567 0 nch W=1.4U L=0.24U
M2 N1N563 E GVSS 0 nch W=1U L=0.24U
M5 N1N567 N1N563 GVSS 0 nch W=1.3U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbh1s5 Q E DIN
M6 N1N565 DIN VDD VDD pch W=4U L=0.24U
M1 N1N563 E VDD VDD pch W=3U L=0.24U
M3 N1N565 E VDD VDD pch W=3.1U L=0.24U
M9 Q N1N565 VDD VDD pch W=6.3U L=0.24U
M7 N1N567 N1N563 N1N565 VDD pch W=4.9U L=0.24U
M8 N1N567 DIN GVSS 0 nch W=1.4U L=0.24U
M10 Q N1N567 GVSS 0 nch W=3.1U L=0.24U
M4 N1N565 E N1N567 0 nch W=3.1U L=0.24U
M2 N1N563 E GVSS 0 nch W=1.8U L=0.24U
M5 N1N567 N1N563 GVSS 0 nch W=1.4U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbh1s6 Q E DIN
M6 N1N565 DIN VDD VDD pch W=4.8U L=0.24U
M1 N1N563 E VDD VDD pch W=3.6U L=0.24U
M3 N1N565 E VDD VDD pch W=3.7U L=0.24U
M9 Q N1N565 VDD VDD pch W=7.6U L=0.24U
M7 N1N567 N1N563 N1N565 VDD pch W=5.9U L=0.24U
M8 N1N567 DIN GVSS 0 nch W=1.8U L=0.24U
M10 Q N1N567 GVSS 0 nch W=3.8U L=0.24U
M4 N1N565 E N1N567 0 nch W=3.7U L=0.24U
M2 N1N563 E GVSS 0 nch W=2.2U L=0.24U
M5 N1N567 N1N563 GVSS 0 nch W=1.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbl1s1 Q EB DIN
M2 N1N260 DIN GVSS 0 nch W=0.9U L=0.24U
M1 N1N260 DIN VDD VDD pch W=1.5U L=0.24U
M4 N1N276 EB GVSS 0 nch W=0.8U L=0.24U
M3 N1N276 EB VDD VDD pch W=1.3U L=0.24U
M8 N1N267 N1N260 GVSS 0 nch W=0.94U L=0.24U
M7 Q N1N276 N1N267 0 nch W=0.94U L=0.24U
M6 Q EB N1N262 VDD pch W=2.6U L=0.24U
M5 N1N262 N1N260 VDD VDD pch W=2.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbl1s2 Q EB DIN
M2 N1N260 DIN GVSS 0 nch W=0.9U L=0.24U
M1 N1N260 DIN VDD VDD pch W=1.6U L=0.24U
M4 N1N276 EB GVSS 0 nch W=0.9U L=0.24U
M3 N1N276 EB VDD VDD pch W=1.8U L=0.24U
M8 N1N267 N1N260 GVSS 0 nch W=1.26U L=0.24U
M7 Q N1N276 N1N267 0 nch W=1.26U L=0.24U
M6 Q EB N1N262 VDD pch W=3.5U L=0.24U
M5 N1N262 N1N260 VDD VDD pch W=3.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbl1s3 Q EB DIN
M4 N1N259 DIN GVSS 0 nch W=1.9U L=0.24U
M2 N1N257 DIN VDD VDD pch W=1.5U L=0.24U
M3 N1N259 EB N1N257 VDD pch W=1.6U L=0.24U
M5 N1N257 N1N285 VDD VDD pch W=1U L=0.24U
M6 N1N257 N1N285 N1N259 0 nch W=1.5U L=0.24U
M7 N1N259 EB GVSS 0 nch W=1U L=0.24U
M9 Q N1N259 GVSS 0 nch W=1.46U L=0.24U
M8 Q N1N257 VDD VDD pch W=2.42U L=0.24U
M1 N1N285 EB VDD VDD pch W=1.3U L=0.24U
M10 N1N285 EB GVSS 0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbl1s4 Q EB DIN
M4 N1N259 DIN GVSS 0 nch W=2.5U L=0.24U
M2 N1N257 DIN VDD VDD pch W=2.8U L=0.24U
M3 N1N259 EB N1N257 VDD pch W=2.8U L=0.24U
M5 N1N257 N1N285 VDD VDD pch W=1.7U L=0.24U
M6 N1N257 N1N285 N1N259 0 nch W=1.8U L=0.24U
M7 N1N259 EB GVSS 0 nch W=1.6U L=0.24U
M9 Q N1N259 GVSS 0 nch W=1.92U L=0.24U
M8 Q N1N257 VDD VDD pch W=4U L=0.24U
M1 N1N285 EB VDD VDD pch W=1.7U L=0.24U
M10 N1N285 EB GVSS 0 nch W=0.9U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbl1s5 Q EB DIN
M4 N1N259 DIN GVSS 0 nch W=3.1U L=0.24U
M2 N1N257 DIN VDD VDD pch W=3.5U L=0.24U
M3 N1N259 EB N1N257 VDD pch W=3.8U L=0.24U
M5 N1N257 N1N285 VDD VDD pch W=2.1U L=0.24U
M6 N1N257 N1N285 N1N259 0 nch W=2.2U L=0.24U
M7 N1N259 EB GVSS 0 nch W=1.6U L=0.24U
M9 Q N1N259 GVSS 0 nch W=3.1U L=0.24U
M8 Q N1N257 VDD VDD pch W=7U L=0.24U
M1 N1N285 EB VDD VDD pch W=2.2U L=0.24U
M10 N1N285 EB GVSS 0 nch W=1U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_tnbl1s6 Q EB DIN
M4 N1N259 DIN GVSS 0 nch W=3.7U L=0.24U
M2 N1N257 DIN VDD VDD pch W=4.2U L=0.24U
M3 N1N259 EB N1N257 VDD pch W=4.6U L=0.24U
M5 N1N257 N1N285 VDD VDD pch W=2.5U L=0.24U
M6 N1N257 N1N285 N1N259 0 nch W=2.6U L=0.24U
M7 N1N259 EB GVSS 0 nch W=1.9U L=0.24U
M9 Q N1N259 GVSS 0 nch W=3.7U L=0.24U
M8 Q N1N257 VDD VDD pch W=8.6U L=0.24U
M1 N1N285 EB VDD VDD pch W=2.6U L=0.24U
M10 N1N285 EB GVSS 0 nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xnr2s1 Q DIN1 DIN2
M9 Q N1N89 VDD VDD pch W=3.1U L=0.24U 
M10 Q N1N89 GVSS 0 nch W=1.1U L=0.24U 
M4 N1N123 DIN1 GVSS 0 nch W=0.6U L=0.24U 
M3 N1N123 DIN1 VDD VDD pch W=1.5U L=0.24U 
M2 N1N83 DIN2 GVSS 0 nch W=0.6U L=0.24U 
M1 N1N83 DIN2 VDD VDD pch W=1.3U L=0.24U 
M5 N1N89 DIN1 DIN2 VDD pch W=1.4U L=0.24U 
M6 DIN2 N1N123 N1N89 0 nch W=0.6U L=0.24U 
M8 N1N83 DIN1 N1N89 0 nch W=0.6U L=0.24U 
M7 N1N89 N1N123 N1N83 VDD pch W=1.4U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xnr2s2 Q DIN1 DIN2
M10 Q N1N89 GVSS 0 nch W=2.2U L=0.24U 
M4 N1N83 DIN1 GVSS 0 nch W=1.2U L=0.24U 
M3 N1N83 DIN1 VDD VDD pch W=3U L=0.24U 
M2 N1N121 DIN2 GVSS 0 nch W=1.5U L=0.24U 
M1 N1N121 DIN2 VDD VDD pch W=2.8U L=0.24U 
M5 N1N89 DIN1 DIN2 VDD pch W=2U L=0.24U 
M6 DIN2 N1N83 N1N89 0 nch W=0.8U L=0.24U 
M8 N1N121 DIN1 N1N89 0 nch W=0.8U L=0.24U 
M7 N1N89 N1N83 N1N121 VDD pch W=2U L=0.24U 
M9 Q N1N89 VDD VDD pch W=5.5U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xnr2s3 Q DIN1 DIN2
M10 Q N1N89 GVSS 0 nch W=3.8U L=0.24U 
M4 N1N83 DIN1 GVSS 0 nch W=2.4U L=0.24U 
M3 N1N83 DIN1 VDD VDD pch W=5.8U L=0.24U 
M2 N1N121 DIN2 GVSS 0 nch W=2.9U L=0.24U 
M1 N1N121 DIN2 VDD VDD pch W=5.2U L=0.24U 
M5 N1N89 DIN1 DIN2 VDD pch W=3U L=0.24U 
M6 DIN2 N1N83 N1N89 0 nch W=1.2U L=0.24U 
M8 N1N121 DIN1 N1N89 0 nch W=1.2U L=0.24U 
M7 N1N89 N1N83 N1N121 VDD pch W=3U L=0.24U 
M9 Q N1N89 VDD VDD pch W=9.5U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xnr3s1 Q DIN1 DIN2 DIN3
M20 Q N1N299 GVSS 0 nch W=2.9U L=0.24U 
M19 Q N1N299 VDD VDD pch W=3.8U L=0.24U 
M15 N1N299 N1N328 DIN2 VDD pch W=1.5U L=0.24U 
M16 DIN2 N1N321 N1N299 0 nch W=0.6U L=0.24U 
M2 N1N309 DIN1 GVSS 0 nch W=1.1U L=0.24U 
M1 N1N309 DIN1 VDD VDD pch W=2.6U L=0.24U 
M4 N1N313 DIN2 GVSS 0 nch W=0.6U L=0.24U 
M3 N1N313 DIN2 VDD VDD pch W=1.8U L=0.24U 
M6 N1N317 DIN3 GVSS 0 nch W=1.2U L=0.24U 
M5 N1N317 DIN3 VDD VDD pch W=2.4U L=0.24U 
M8 N1N317 N1N309 N1N321 0 nch W=0.7U L=0.24U 
M7 N1N321 DIN1 N1N317 VDD pch W=1.7U L=0.24U 
M10 DIN3 DIN1 N1N321 0 nch W=0.7U L=0.24U 
M9 N1N321 N1N309 DIN3 VDD pch W=1.7U L=0.24U 
M11 N1N328 DIN1 DIN3 VDD pch W=1.7U L=0.24U 
M12 DIN3 N1N309 N1N328 0 nch W=0.7U L=0.24U 
M13 N1N328 N1N309 N1N317 VDD pch W=1.7U L=0.24U 
M14 N1N317 DIN1 N1N328 0 nch W=0.7U L=0.24U 
M18 N1N313 N1N328 N1N299 0 nch W=0.6U L=0.24U 
M17 N1N299 N1N321 N1N313 VDD pch W=1.5U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xnr3s2 Q DIN1 DIN2 DIN3
M20 Q N1N299 GVSS 0 nch W=4.4U L=0.24U 
M19 Q N1N299 VDD VDD pch W=5.7U L=0.24U 
M15 N1N299 N1N328 DIN2 VDD pch W=2.1U L=0.24U 
M16 DIN2 N1N321 N1N299 0 nch W=0.8U L=0.24U 
M2 N1N309 DIN1 GVSS 0 nch W=1.7U L=0.24U 
M1 N1N309 DIN1 VDD VDD pch W=3.9U L=0.24U 
M4 N1N313 DIN2 GVSS 0 nch W=1U L=0.24U 
M3 N1N313 DIN2 VDD VDD pch W=2.6U L=0.24U 
M6 N1N317 DIN3 GVSS 0 nch W=1.8U L=0.24U 
M5 N1N317 DIN3 VDD VDD pch W=3.6U L=0.24U 
M8 N1N317 N1N309 N1N321 0 nch W=1U L=0.24U 
M7 N1N321 DIN1 N1N317 VDD pch W=2.4U L=0.24U 
M10 DIN3 DIN1 N1N321 0 nch W=1U L=0.24U 
M9 N1N321 N1N309 DIN3 VDD pch W=2.4U L=0.24U 
M11 N1N328 DIN1 DIN3 VDD pch W=2.4U L=0.24U 
M12 DIN3 N1N309 N1N328 0 nch W=1U L=0.24U 
M13 N1N328 N1N309 N1N317 VDD pch W=2.4U L=0.24U 
M14 N1N317 DIN1 N1N328 0 nch W=1U L=0.24U 
M18 N1N313 N1N328 N1N299 0 nch W=0.8U L=0.24U 
M17 N1N299 N1N321 N1N313 VDD pch W=2.1U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xnr3s3 Q DIN1 DIN2 DIN3
M20 Q N1N299 GVSS 0 nch W=7.1U L=0.24U 
M19 Q N1N299 VDD VDD pch W=9.5U L=0.24U 
M15 N1N299 N1N328 DIN2 VDD pch W=3.2U L=0.24U 
M16 DIN2 N1N321 N1N299 0 nch W=1.2U L=0.24U 
M2 N1N309 DIN1 GVSS 0 nch W=3.1U L=0.24U 
M1 N1N309 DIN1 VDD VDD pch W=7U L=0.24U 
M4 N1N313 DIN2 GVSS 0 nch W=1.8U L=0.24U 
M3 N1N313 DIN2 VDD VDD pch W=4.4U L=0.24U 
M6 N1N317 DIN3 GVSS 0 nch W=3.2U L=0.24U 
M5 N1N317 DIN3 VDD VDD pch W=6.5U L=0.24U 
M8 N1N317 N1N309 N1N321 0 nch W=1.5U L=0.24U 
M7 N1N321 DIN1 N1N317 VDD pch W=3.6U L=0.24U 
M10 DIN3 DIN1 N1N321 0 nch W=1.5U L=0.24U 
M9 N1N321 N1N309 DIN3 VDD pch W=3.6U L=0.24U 
M11 N1N328 DIN1 DIN3 VDD pch W=3.6U L=0.24U 
M12 DIN3 N1N309 N1N328 0 nch W=1.5U L=0.24U 
M13 N1N328 N1N309 N1N317 VDD pch W=3.6U L=0.24U 
M14 N1N317 DIN1 N1N328 0 nch W=1.5U L=0.24U 
M18 N1N313 N1N328 N1N299 0 nch W=1.2U L=0.24U 
M17 N1N299 N1N321 N1N313 VDD pch W=3.2U L=0.24U 
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xor2s1 Q DIN1 DIN2
M2       N1N83 DIN1 GVSS    0 nch W=0.6U L=0.24U
M1       N1N83 DIN1 VDD  VDD pch W=1.3U L=0.24U
M4       N1N85 DIN2 GVSS    0 nch W=0.6U L=0.24U
M3       N1N85 DIN2 VDD  VDD pch W=1.5U L=0.24U
M5       N1N91 DIN2 N1N83  VDD pch W=1.4U L=0.24U
M6       N1N83 N1N85 N1N91  0 nch W=0.6U L=0.24U
M8       DIN1 DIN2 N1N91  0 nch W=0.6U L=0.24U
M7       N1N91 N1N85 DIN1  VDD pch W=1.4U L=0.24U
M10      Q N1N91 GVSS    0 nch W=1.9U L=0.24U
M9       Q N1N91 VDD  VDD pch W=2.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xor2s2 Q DIN1 DIN2
M2       N1N83 DIN1 GVSS    0 nch W=1.2U L=0.24U
M1       N1N83 DIN1 VDD  VDD pch W=2.6U L=0.24U
M4       N1N85 DIN2 GVSS    0 nch W=1.2U L=0.24U
M3       N1N85 DIN2 VDD  VDD pch W=3.0U L=0.24U
M5       N1N91 DIN2 N1N83  VDD pch W=2.0U L=0.24U
M6       N1N83 N1N85 N1N91  0 nch W=0.8U L=0.24U
M8       DIN1 DIN2 N1N91  0 nch W=0.8U L=0.24U
M7       N1N91 N1N85 DIN1  VDD pch W=2.0U L=0.24U
M10      Q N1N91 GVSS    0 nch W=3.7U L=0.24U
M9       Q N1N91 VDD  VDD pch W=5.0U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xor2s3 Q DIN1 DIN2
M2       N1N83 DIN1 GVSS    0 nch W=2.4U L=0.24U
M1       N1N83 DIN1 VDD  VDD pch W=5.2U L=0.24U
M4       N1N85 DIN2 GVSS    0 nch W=2.4U L=0.24U
M3       N1N85 DIN2 VDD  VDD pch W=5.8U L=0.24U
M5       N1N91 DIN2 N1N83  VDD pch W=3.0U L=0.24U
M6       N1N83 N1N85 N1N91  0 nch W=1.2U L=0.24U
M8       DIN1 DIN2 N1N91  0 nch W=1.2U L=0.24U
M7       N1N91 N1N85 DIN1  VDD pch W=3.0U L=0.24U
M10      Q N1N91 GVSS    0 nch W=6.7U L=0.24U
M9       Q N1N91 VDD  VDD pch W=9.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xor3s1 Q DIN1 DIN2 DIN3
M20      Q N1N307 GVSS    0 nch W=2.9U L=0.24U
M19      Q N1N307 VDD  VDD pch W=3.8U L=0.24U
M15      N1N307 DIN2 N1N311  VDD pch W=1.5U L=0.24U
M16      N1N311 N1N321 N1N307  0 nch W=0.6U L=0.24U
M2       N1N360 DIN1 GVSS    0 nch W=1.1U L=0.24U
M1       N1N360 DIN1 VDD  VDD pch W=2.6U L=0.24U
M4       N1N321 DIN2 GVSS    0 nch W=0.7U L=0.24U
M3       N1N321 DIN2 VDD  VDD pch W=1.4U L=0.24U
M6       N1N325 DIN3 GVSS    0 nch W=1.2U L=0.24U
M5       N1N325 DIN3 VDD  VDD pch W=2.4U L=0.24U
M7       N1N311 DIN1 N1N325  VDD pch W=1.7U L=0.24U
M8       N1N325 N1N360 N1N311  0 nch W=0.7U L=0.24U
M10      DIN3 DIN1 N1N311  0 nch W=0.7U L=0.24U
M9       N1N311 N1N360 DIN3  VDD pch W=1.7U L=0.24U
M12      DIN3 N1N360 N1N338  0 nch W=0.7U L=0.24U
M11      N1N338 DIN1 DIN3  VDD pch W=1.7U L=0.24U
M13      N1N338 N1N360 N1N325  VDD pch W=1.7U L=0.24U
M14      N1N325 DIN1 N1N338  0 nch W=0.7U L=0.24U
M17      N1N307 N1N321 N1N338  VDD pch W=1.5U L=0.24U
M18      N1N338 DIN2 N1N307  0 nch W=0.6U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xor3s2 Q DIN1 DIN2 DIN3
M20      Q N1N307 GVSS    0 nch W=4.4U L=0.24U
M19      Q N1N307 VDD  VDD pch W=5.7U L=0.24U
M15      N1N307 DIN2 N1N311  VDD pch W=2.1U L=0.24U
M16      N1N311 N1N321 N1N307  0 nch W=0.8U L=0.24U
M2       N1N360 DIN1 GVSS    0 nch W=1.7U L=0.24U
M1       N1N360 DIN1 VDD  VDD pch W=3.9U L=0.24U
M4       N1N321 DIN2 GVSS    0 nch W=1.1U L=0.24U
M3       N1N321 DIN2 VDD  VDD pch W=2.1U L=0.24U
M6       N1N325 DIN3 GVSS    0 nch W=1.8U L=0.24U
M5       N1N325 DIN3 VDD  VDD pch W=3.6U L=0.24U
M7       N1N311 DIN1 N1N325  VDD pch W=2.4U L=0.24U
M8       N1N325 N1N360 N1N311  0 nch W=1.0U L=0.24U
M10      DIN3 DIN1 N1N311  0 nch W=1.0U L=0.24U
M9       N1N311 N1N360 DIN3  VDD pch W=2.4U L=0.24U
M12      DIN3 N1N360 N1N338  0 nch W=1.0U L=0.24U
M11      N1N338 DIN1 DIN3  VDD pch W=2.4U L=0.24U
M13      N1N338 N1N360 N1N325  VDD pch W=2.4U L=0.24U
M14      N1N325 DIN1 N1N338  0 nch W=1.0U L=0.24U
M17      N1N307 N1N321 N1N338  VDD pch W=2.1U L=0.24U
M18      N1N338 DIN2 N1N307  0 nch W=0.8U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_xor3s3 Q DIN1 DIN2 DIN3
M20      Q N1N307 GVSS    0 nch W=7.1U L=0.24U
M19      Q N1N307 VDD  VDD pch W=9.54U L=0.24U
M15      N1N307 DIN2 N1N311  VDD pch W=3.2U L=0.24U
M16      N1N311 N1N321 N1N307  0 nch W=1.2U L=0.24U
M2       N1N360 DIN1 GVSS    0 nch W=3.1U L=0.24U
M1       N1N360 DIN1 VDD  VDD pch W=7.0U L=0.24U
M4       N1N321 DIN2 GVSS    0 nch W=2.0U L=0.24U
M3       N1N321 DIN2 VDD  VDD pch W=3.8U L=0.24U
M6       N1N325 DIN3 GVSS    0 nch W=3.2U L=0.24U
M5       N1N325 DIN3 VDD  VDD pch W=6.5U L=0.24U
M7       N1N311 DIN1 N1N325  VDD pch W=3.6U L=0.24U
M8       N1N325 N1N360 N1N311  0 nch W=1.5U L=0.24U
M10      DIN3 DIN1 N1N311  0 nch W=1.5U L=0.24U
M9       N1N311 N1N360 DIN3  VDD pch W=3.6U L=0.24U
M12      DIN3 N1N360 N1N338  0 nch W=1.5U L=0.24U
M11      N1N338 DIN1 DIN3  VDD pch W=3.6U L=0.24U
M13      N1N338 N1N360 N1N325  VDD pch W=3.6U L=0.24U
M14      N1N325 DIN1 N1N338  0 nch W=1.5U L=0.24U
M17      N1N307 N1N321 N1N338  VDD pch W=3.2U L=0.24U
M18      N1N338 DIN2 N1N307  0 nch W=1.2U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_avdd PAD AVDD
C1I4110 PAD N1I41TP0 235FF
C1I4111 N1I41TP2 PAD 235FF
M1 AVDD N1N17 AVSS AVSS nch W=300U L=0.34U
M1I410 N1I41TP7 N1I41TP0 NVDD NVDD pch W=38U L=0.34U
M1I411 N1I41TP0 N1I41TP1 NVDD NVDD pch W=6U L=6U
M1I412 N1I41TP2 N1I41TP3 NVSS NVSS nch W=6U L=6U
M1I413 N1I41TP4 N1I41TP2 N1I41TP5 NVSS nch W=38U L=0.34U
R1 N1N17 AVSS 400
R1I414 N1I41TP7 EVSS 123
R1I415 NVDD N1I41TP3 198
R1I416 EVDD N1I41TP4 177
R1I417 N1I41TP1 NVSS 198
R1I418 N1I41TP5 NVSS 0.21
R1I419 N1I41TP5 NVSS 0.21
R2 AVDD PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_avss PAD AVSS
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 AVSS N1N48 AVDD AVDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 AVDD N1N48 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 AVSS PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cainr25s4 PAD Q
C1I35710 PAD N1I357TP0 235FF
C1I35711 N1I357TP2 PAD 235FF
M1I3570 N1I357TP7 N1I357TP0 NVDD NVDD pch W=38U L=0.34U
M1I3571 N1I357TP0 N1I357TP1 NVDD NVDD pch W=6U L=6U
M1I3572 N1I357TP2 N1I357TP3 NVSS NVSS nch W=6U L=6U
M1I3573 N1I357TP4 N1I357TP2 N1I357TP5 NVSS nch W=38U L=0.34U
R1 PAD Q 200
R1I3574 N1I357TP7 EVSS 123
R1I3575 NVDD N1I357TP3 198
R1I3576 EVDD N1I357TP4 177
R1I3577 N1I357TP1 NVSS 198
R1I3578 N1I357TP5 NVSS 0.21
R1I3579 N1I357TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_caon25s4 PAD DIN
C1I36910 PAD N1I369TP0 235FF
C1I36911 N1I369TP2 PAD 235FF
M1I3690 N1I369TP7 N1I369TP0 NVDD NVDD pch W=38U L=0.34U
M1I3691 N1I369TP0 N1I369TP1 NVDD NVDD pch W=6U L=6U
M1I3692 N1I369TP2 N1I369TP3 NVSS NVSS nch W=6U L=6U
M1I3693 N1I369TP4 N1I369TP2 N1I369TP5 NVSS nch W=38U L=0.34U
R1 PAD DIN 0.30
R1I3694 N1I369TP7 EVSS 123
R1I3695 NVDD N1I369TP3 198
R1I3696 EVDD N1I369TP4 177
R1I3697 N1I369TP1 NVSS 198
R1I3698 N1I369TP5 NVSS 0.21
R1I3699 N1I369TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cdavdd AVDD PAD VDD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 VDD N1N17 GVSS 0 nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N17 GVSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 VDD PAD 0.002
R3 AVDD VDD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cdavss AVSS PAD VSS
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 GVSS N1N48 VDD VDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 VDD N1N48 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 GVSS PAD 0.002
R3 AVSS GVSS 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cdvdd PAD VDD N1
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 VDD N1N17 GVSS 0 nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N17 GVSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 VDD PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cdvss PAD GVSS N1
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 GVSS N1N48 VDD VDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 VDD N1N48 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 GVSS PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cii25s1 PAD Q
C1I38610 PAD N1I386TP0 235FF
C1I38611 N1I386TP2 PAD 235FF
M1 Q TP2 VDD VDD pch W=3.8U L=0.24U
M1I3860 N1I386TP7 N1I386TP0 NVDD NVDD pch W=38U L=0.34U
M1I3861 N1I386TP0 N1I386TP1 NVDD NVDD pch W=6U L=6U
M1I3862 N1I386TP2 N1I386TP3 NVSS NVSS nch W=6U L=6U
M1I3863 N1I386TP4 N1I386TP2 N1I386TP5 NVSS nch W=38U L=0.34U
M2 Q TP2 GVSS 0 nch W=1.36U L=0.24U
M6 TP2 VDD VDD VDD pch W=100U L=0.48U
M7 TP2 GVSS VSS 0 nch W=100U L=0.48U
R1 TP2 PAD 300
R1I3864 N1I386TP7 EVSS 123
R1I3865 NVDD N1I386TP3 198
R1I3866 EVDD N1I386TP4 177
R1I3867 N1I386TP1 NVSS 198
R1I3868 N1I386TP5 NVSS 0.21
R1I3869 N1I386TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cii25s4 PAD Q
C1I39610 PAD N1I396TP0 235FF
C1I39611 N1I396TP2 PAD 235FF
M1 Q TP2 VDD VDD pch W=30U L=0.24U
M1I3960 N1I396TP7 N1I396TP0 NVDD NVDD pch W=38U L=0.34U
M1I3961 N1I396TP0 N1I396TP1 NVDD NVDD pch W=6U L=6U
M1I3962 N1I396TP2 N1I396TP3 NVSS NVSS nch W=6U L=6U
M1I3963 N1I396TP4 N1I396TP2 N1I396TP5 NVSS nch W=38U L=0.34U
M2 Q TP2 GVSS 0 nch W=10.12U L=0.24U
M6 TP2 VDD VDD VDD pch W=100U L=0.48U
M7 TP2 GVSS VSS 0 nch W=100U L=0.48U
R1 TP2 PAD 300
R1I3964 N1I396TP7 EVSS 123
R1I3965 NVDD N1I396TP3 198
R1I3966 EVDD N1I396TP4 177
R1I3967 N1I396TP1 NVSS 198
R1I3968 N1I396TP5 NVSS 0.21
R1I3969 N1I396TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ciis25s1 PAD Q
C1I50810 PAD N1I508TP0 235FF
C1I50811 N1I508TP2 PAD 235FF
M1 TP0 TP5 VDD VDD pch W=2.74U L=0.24U
M1I5080 N1I508TP7 N1I508TP0 NVDD NVDD pch W=38U L=0.34U
M1I5081 N1I508TP0 N1I508TP1 NVDD NVDD pch W=6U L=6U
M1I5082 N1I508TP2 N1I508TP3 NVSS NVSS nch W=6U L=6U
M1I5083 N1I508TP4 N1I508TP2 N1I508TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP5 TP0 VDD pch W=2.74U L=0.24U
M3 TP1 TP5 TP2 0 nch W=24U L=0.24U
M4 TP2 TP5 GVSS 0 nch W=24U L=0.24U
M5 GVSS TP1 TP0 VDD pch W=7.8U L=0.24U
M6 TP2 TP1 VDD 0 nch W=0.4U L=0.24U
M7 TP3 TP1 VDD VDD pch W=1U L=0.24U
M8 TP3 TP1 GVSS 0 nch W=8.2U L=0.24U
M9 Q TP3 VDD VDD pch W=17.5U L=0.24U
M10 Q TP3 GVSS 0 nch W=1U L=0.24U
M13 TP5 VDD VDD VDD pch W=100U L=0.48U
M14 TP5 GVSS VSS 0 nch W=100U L=0.48U
R1 PAD TP5 300
R1I5084 N1I508TP7 EVSS 123
R1I5085 NVDD N1I508TP3 198
R1I5086 EVDD N1I508TP4 177
R1I5087 N1I508TP1 NVSS 198
R1I5088 N1I508TP5 NVSS 0.21
R1I5089 N1I508TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ciis25s4 PAD Q
C1I49710 PAD N1I497TP0 235FF
C1I49711 N1I497TP2 PAD 235FF
M1 TP0 TP5 VDD VDD pch W=2.74U L=0.24U
M1I4970 N1I497TP7 N1I497TP0 NVDD NVDD pch W=38U L=0.34U
M1I4971 N1I497TP0 N1I497TP1 NVDD NVDD pch W=6U L=6U
M1I4972 N1I497TP2 N1I497TP3 NVSS NVSS nch W=6U L=6U
M1I4973 N1I497TP4 N1I497TP2 N1I497TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP5 TP0 VDD pch W=2.74U L=0.24U
M3 TP1 TP5 TP2 0 nch W=42U L=0.24U
M4 TP2 TP5 GVSS 0 nch W=42U L=0.24U
M5 GVSS TP1 TP0 VDD pch W=4.8U L=0.24U
M6 TP2 TP1 VDD 0 nch W=0.4U L=0.24U
M7 TP3 TP1 VDD VDD pch W=1U L=0.24U
M8 TP3 TP1 GVSS 0 nch W=8.5U L=0.24U
M9 Q TP3 VDD VDD pch W=15.2U L=0.24U
M10 Q TP3 GVSS 0 nch W=1.1U L=0.24U
M13 TP5 VDD VDD VDD pch W=100U L=0.48U
M14 TP5 GVSS VSS 0 nch W=100U L=0.48U
R1 PAD TP5 300
R1I4974 N1I497TP7 EVSS 123
R1I4975 NVDD N1I497TP3 198
R1I4976 EVDD N1I497TP4 177
R1I4977 N1I497TP1 NVSS 198
R1I4978 N1I497TP5 NVSS 0.21
R1I4979 N1I497TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cin25s1 PAD Q
C1I38610 PAD N1I386TP0 235FF
C1I38611 N1I386TP2 PAD 235FF
M1 TP1 TP2 VDD VDD pch W=3.8U L=0.24U
M1I3860 N1I386TP7 N1I386TP0 NVDD NVDD pch W=38U L=0.34U
M1I3861 N1I386TP0 N1I386TP1 NVDD NVDD pch W=6U L=6U
M1I3862 N1I386TP2 N1I386TP3 NVSS NVSS nch W=6U L=6U
M1I3863 N1I386TP4 N1I386TP2 N1I386TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP2 GVSS 0 nch W=1.36U L=0.24U
M3 Q TP1 VDD VDD pch W=5.6U L=0.24U
M4 Q TP1 GVSS 0 nch W=2.6U L=0.24U
M6 TP2 VDD VDD VDD pch W=100U L=0.48U
M7 TP2 GVSS VSS 0 nch W=100U L=0.48U
R1 TP2 PAD 300
R1I3864 N1I386TP7 EVSS 123
R1I3865 NVDD N1I386TP3 198
R1I3866 EVDD N1I386TP4 177
R1I3867 N1I386TP1 NVSS 198
R1I3868 N1I386TP5 NVSS 0.21
R1I3869 N1I386TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cin25s4 PAD Q
C1I39610 PAD N1I396TP0 235FF
C1I39611 N1I396TP2 PAD 235FF
M1 TP1 TP2 VDD VDD pch W=30U L=0.24U
M1I3960 N1I396TP7 N1I396TP0 NVDD NVDD pch W=38U L=0.34U
M1I3961 N1I396TP0 N1I396TP1 NVDD NVDD pch W=6U L=6U
M1I3962 N1I396TP2 N1I396TP3 NVSS NVSS nch W=6U L=6U
M1I3963 N1I396TP4 N1I396TP2 N1I396TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP2 GVSS 0 nch W=10.12U L=0.24U
M3 Q TP1 VDD VDD pch W=35.52U L=0.24U
M4 Q TP1 GVSS 0 nch W=15.92U L=0.24U
M6 TP2 VDD VDD VDD pch W=100U L=0.48U
M7 TP2 GVSS VSS 0 nch W=100U L=0.48U
R1 TP2 PAD 300
R1I3964 N1I396TP7 EVSS 123
R1I3965 NVDD N1I396TP3 198
R1I3966 EVDD N1I396TP4 177
R1I3967 N1I396TP1 NVSS 198
R1I3968 N1I396TP5 NVSS 0.21
R1I3969 N1I396TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cins25s1 PAD Q
C1I50810 PAD N1I508TP0 235FF
C1I50811 N1I508TP2 PAD 235FF
M1 TP0 TP5 VDD VDD pch W=2.74U L=0.24U
M1I5080 N1I508TP7 N1I508TP0 NVDD NVDD pch W=38U L=0.34U
M1I5081 N1I508TP0 N1I508TP1 NVDD NVDD pch W=6U L=6U
M1I5082 N1I508TP2 N1I508TP3 NVSS NVSS nch W=6U L=6U
M1I5083 N1I508TP4 N1I508TP2 N1I508TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP5 TP0 VDD pch W=2.74U L=0.24U
M3 TP1 TP5 TP2 0 nch W=24U L=0.24U
M4 TP2 TP5 GVSS 0 nch W=24U L=0.24U
M5 GVSS TP1 TP0 VDD pch W=7.8U L=0.24U
M6 TP2 TP1 VDD 0 nch W=0.4U L=0.24U
M7 TP3 TP1 VDD VDD pch W=1U L=0.24U
M8 TP3 TP1 GVSS 0 nch W=8.2U L=0.24U
M9 TP4 TP3 VDD VDD pch W=17.5U L=0.24U
M10 TP4 TP3 GVSS 0 nch W=1U L=0.24U
M11 Q TP4 VDD VDD pch W=8.2U L=0.24U
M12 Q TP4 GVSS 0 nch W=4.1U L=0.24U
M13 TP5 VDD VDD VDD pch W=100U L=0.48U
M14 TP5 GVSS VSS 0 nch W=100U L=0.48U
R1 PAD TP5 300
R1I5084 N1I508TP7 EVSS 123
R1I5085 NVDD N1I508TP3 198
R1I5086 EVDD N1I508TP4 177
R1I5087 N1I508TP1 NVSS 198
R1I5088 N1I508TP5 NVSS 0.21
R1I5089 N1I508TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cins25s4 PAD Q
C1I49510 PAD N1I495TP0 235FF
C1I49511 N1I495TP2 PAD 235FF
M1 TP0 TP5 VDD VDD pch W=2.74U L=0.24U
M1I4950 N1I495TP7 N1I495TP0 NVDD NVDD pch W=38U L=0.34U
M1I4951 N1I495TP0 N1I495TP1 NVDD NVDD pch W=6U L=6U
M1I4952 N1I495TP2 N1I495TP3 NVSS NVSS nch W=6U L=6U
M1I4953 N1I495TP4 N1I495TP2 N1I495TP5 NVSS nch W=38U L=0.34U
M2 TP1 TP5 TP0 VDD pch W=2.74U L=0.24U
M3 TP1 TP5 TP2 0 nch W=42U L=0.24U
M4 TP2 TP5 GVSS 0 nch W=42U L=0.24U
M5 GVSS TP1 TP0 VDD pch W=4.8U L=0.24U
M6 TP2 TP1 VDD 0 nch W=0.4U L=0.24U
M7 TP3 TP1 VDD VDD pch W=1U L=0.24U
M8 TP3 TP1 GVSS 0 nch W=8.5U L=0.24U
M9 TP4 TP3 VDD VDD pch W=15.2U L=0.24U
M10 TP4 TP3 GVSS 0 nch W=1.1U L=0.24U
M11 Q TP4 VDD VDD pch W=30.1U L=0.24U
M12 Q TP4 GVSS 0 nch W=18.5U L=0.24U
M13 TP5 VDD VDD VDD pch W=100U L=0.48U
M14 TP5 GVSS VSS 0 nch W=100U L=0.48U
R1 PAD TP5 300
R1I4954 N1I495TP7 EVSS 123
R1I4955 NVDD N1I495TP3 198
R1I4956 EVDD N1I495TP4 177
R1I4957 N1I495TP1 NVSS 198
R1I4958 N1I495TP5 NVSS 0.21
R1I4959 N1I495TP5 NVSS 0.21
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cioit25s1 DIN E PAD Q
C1I35310 PAD N1I353TP0 235FF
C1I35311 N1I353TP2 PAD 235FF
M1I3530 N1I353TP7 N1I353TP0 NVDD NVDD pch W=38U L=0.34U
M1I3531 N1I353TP0 N1I353TP1 NVDD NVDD pch W=6U L=6U
M1I3532 N1I353TP2 N1I353TP3 NVSS NVSS nch W=6U L=6U
M1I3533 N1I353TP4 N1I353TP2 N1I353TP5 NVSS nch W=38U L=0.34U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E GVSS 0 nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=13U L=0.24U
M6 TP2 E TP3 0 nch W=10U L=0.24U
M7 TP3 TP1 GVSS 0 nch W=7U L=0.24U
M8 VDD TP20 TP2 VDD pch W=13U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 GVSS TP20 TP3 0 nch W=7U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=15.5U L=0.34U
M14 TP14 TP3 NVSS 0 nch W=5U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=15.5U L=0.34U
M18 TP15 TP3 NVSS 0 nch W=5U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=15.5U L=0.34U
M22 TP16 TP3 NVSS 0 nch W=5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=15.5U L=0.34U
M26 TP17 TP3 NVSS 0 nch W=5U L=0.34U
M27 PAD NVSS NVSS 0 nch W=34U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 GVSS TP4 Q 0 nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 GVSS TP13 TP4 0 nch W=4.1U L=0.24U
M33 TP20 DIN VDD VDD pch W=5.4U L=0.24U
M34 TP20 DIN GVSS 0 nch W=7U L=0.24U
R1I3534 N1I353TP7 EVSS 123
R1I3535 NVDD N1I353TP3 198
R1I3536 EVDD N1I353TP4 177
R1I3537 N1I353TP1 NVSS 198
R1I3538 N1I353TP5 NVSS 0.21
R1I3539 N1I353TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cioit25s2 DIN E PAD Q
C1I32310 PAD N1I323TP0 235FF
C1I32311 N1I323TP2 PAD 235FF
M1I3230 N1I323TP7 N1I323TP0 NVDD NVDD pch W=38U L=0.34U
M1I3231 N1I323TP0 N1I323TP1 NVDD NVDD pch W=6U L=6U
M1I3232 N1I323TP2 N1I323TP3 NVSS NVSS nch W=6U L=6U
M1I3233 N1I323TP4 N1I323TP2 N1I323TP5 NVSS nch W=38U L=0.34U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E GVSS 0 nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=13U L=0.24U
M6 TP2 E TP3 0 nch W=10U L=0.24U
M7 TP3 TP1 GVSS 0 nch W=7.2U L=0.24U
M8 VDD TP20 TP2 VDD pch W=13U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 GVSS TP20 TP3 0 nch W=7.2U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=35.5U L=0.34U
M14 TP14 TP3 NVSS 0 nch W=10.8U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=35.5U L=0.34U
M18 TP15 TP3 NVSS 0 nch W=10.8U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=35.5U L=0.34U
M22 TP16 TP3 NVSS 0 nch W=10.8U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=35.5U L=0.34U
M26 TP17 TP3 NVSS 0 nch W=10.8U L=0.34U
M27 PAD NVSS NVSS 0 nch W=24U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 GVSS TP4 Q 0 nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 GVSS TP13 TP4 0 nch W=4.1U L=0.24U
M33 TP20 DIN VDD VDD pch W=3U L=0.24U
M34 TP20 DIN GVSS 0 nch W=7U L=0.24U
R1I3234 N1I323TP7 EVSS 123
R1I3235 NVDD N1I323TP3 198
R1I3236 EVDD N1I323TP4 177
R1I3237 N1I323TP1 NVSS 198
R1I3238 N1I323TP5 NVSS 0.21
R1I3239 N1I323TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cioit25s3 DIN E PAD Q
C1I32810 PAD N1I328TP0 235FF
C1I32811 N1I328TP2 PAD 235FF
M1I3280 N1I328TP7 N1I328TP0 NVDD NVDD pch W=38U L=0.34U
M1I3281 N1I328TP0 N1I328TP1 NVDD NVDD pch W=6U L=6U
M1I3282 N1I328TP2 N1I328TP3 NVSS NVSS nch W=6U L=6U
M1I3283 N1I328TP4 N1I328TP2 N1I328TP5 NVSS nch W=38U L=0.34U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E GVSS 0 nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=14U L=0.24U
M6 TP2 E TP3 0 nch W=10U L=0.24U
M7 TP3 TP1 GVSS 0 nch W=7.6U L=0.24U
M8 VDD TP20 TP2 VDD pch W=14U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 GVSS TP20 TP3 0 nch W=7.6U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=84U L=0.34U
M14 TP14 TP3 NVSS 0 nch W=24.5U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=84U L=0.34U
M18 TP15 TP3 NVSS 0 nch W=24.5U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=84U L=0.34U
M22 TP16 TP3 NVSS 0 nch W=24.5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=84U L=0.34U
M26 TP17 TP3 NVSS 0 nch W=24.5U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 GVSS TP4 Q 0 nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 GVSS TP13 TP4 0 nch W=4.1U L=0.24U
M33 TP20 DIN VDD VDD pch W=3U L=0.24U
M34 TP20 DIN GVSS 0 nch W=7U L=0.24U
R1I3284 N1I328TP7 EVSS 123
R1I3285 NVDD N1I328TP3 198
R1I3286 EVDD N1I328TP4 177
R1I3287 N1I328TP1 NVSS 198
R1I3288 N1I328TP5 NVSS 0.21
R1I3289 N1I328TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_cioit25s4 DIN E PAD Q
C1I32410 PAD N1I324TP0 235FF
C1I32411 N1I324TP2 PAD 235FF
M1I3240 N1I324TP7 N1I324TP0 NVDD NVDD pch W=38U L=0.34U
M1I3241 N1I324TP0 N1I324TP1 NVDD NVDD pch W=6U L=6U
M1I3242 N1I324TP2 N1I324TP3 NVSS NVSS nch W=6U L=6U
M1I3243 N1I324TP4 N1I324TP2 N1I324TP5 NVSS nch W=38U L=0.34U
M3 TP20 E VDD VDD pch W=6U L=0.24U
M4 TP20 E GVSS 0 nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=18U L=0.24U
M6 TP2 E TP3 0 nch W=10U L=0.24U
M7 TP3 TP20 GVSS 0 nch W=10U L=0.24U
M8 VDD TP1 TP2 VDD pch W=18U L=0.24U
M9 TP2 TP20 TP3 VDD pch W=10U L=0.24U
M10 GVSS TP1 TP3 0 nch W=10U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=152U L=0.34U
M14 TP14 TP3 NVSS 0 nch W=40.8U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=152U L=0.34U
M18 TP15 TP3 NVSS 0 nch W=40.8U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=152U L=0.34U
M22 TP16 TP3 NVSS 0 nch W=40.5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=152U L=0.34U
M26 TP17 TP3 NVSS 0 nch W=40.8U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 GVSS TP4 Q 0 nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 GVSS TP13 TP4 0 nch W=4.1U L=0.24U
M33 TP1 DIN VDD VDD pch W=3U L=0.24U
M34 TP1 DIN GVSS 0 nch W=7U L=0.24U
R1I3244 N1I324TP7 EVSS 123
R1I3245 NVDD N1I324TP3 198
R1I3246 EVDD N1I324TP4 177
R1I3247 N1I324TP1 NVSS 198
R1I3248 N1I324TP5 NVSS 0.21
R1I3249 N1I324TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ciont25s1 DIN E PAD Q
C1I35310 PAD N1I353TP0 235FF
C1I35311 N1I353TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6U L=0.24U
M1I3530 N1I353TP7 N1I353TP0 NVDD NVDD pch W=38U L=0.34U
M1I3531 N1I353TP0 N1I353TP1 NVDD NVDD pch W=6U L=6U
M1I3532 N1I353TP2 N1I353TP3 NVSS NVSS nch W=6U L=6U
M1I3533 N1I353TP4 N1I353TP2 N1I353TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN GVSS 0 nch W=2U L=0.24U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E GVSS 0 nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=13U L=0.24U
M6 TP2 E TP3 0 nch W=10U L=0.24U
M7 TP3 TP1 GVSS 0 nch W=7U L=0.24U
M8 VDD TP20 TP2 VDD pch W=13U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 GVSS TP20 TP3 0 nch W=7U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=15.5U L=0.34U
M14 TP14 TP3 NVSS 0 nch W=5U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=15.5U L=0.34U
M18 TP15 TP3 NVSS 0 nch W=5U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=15.5U L=0.34U
M22 TP16 TP3 NVSS 0 nch W=5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=15.5U L=0.34U
M26 TP17 TP3 NVSS 0 nch W=5U L=0.34U
M27 PAD NVSS NVSS 0 nch W=34U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 GVSS TP4 Q 0 nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 GVSS TP13 TP4 0 nch W=4.1U L=0.24U
M33 TP20 TP0 VDD VDD pch W=5.4U L=0.24U
M34 TP20 TP0 GVSS 0 nch W=7U L=0.24U
R1I3534 N1I353TP7 EVSS 123
R1I3535 NVDD N1I353TP3 198
R1I3536 EVDD N1I353TP4 177
R1I3537 N1I353TP1 NVSS 198
R1I3538 N1I353TP5 NVSS 0.21
R1I3539 N1I353TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ciont25s2 DIN E PAD Q
C1I32310 PAD N1I323TP0 235FF
C1I32311 N1I323TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6U L=0.24U
M1I3230 N1I323TP7 N1I323TP0 NVDD NVDD pch W=38U L=0.34U
M1I3231 N1I323TP0 N1I323TP1 NVDD NVDD pch W=6U L=6U
M1I3232 N1I323TP2 N1I323TP3 NVSS NVSS nch W=6U L=6U
M1I3233 N1I323TP4 N1I323TP2 N1I323TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN GVSS 0 nch W=2U L=0.24U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E GVSS 0 nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=13U L=0.24U
M6 TP2 E TP3 0 nch W=10U L=0.24U
M7 TP3 TP1 GVSS 0 nch W=7.2U L=0.24U
M8 VDD TP20 TP2 VDD pch W=13U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 GVSS TP20 TP3 0 nch W=7.2U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=35.5U L=0.34U
M14 TP14 TP3 NVSS 0 nch W=10.8U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=35.5U L=0.34U
M18 TP15 TP3 NVSS 0 nch W=10.8U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=35.5U L=0.34U
M22 TP16 TP3 NVSS 0 nch W=10.8U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=35.5U L=0.34U
M26 TP17 TP3 NVSS 0 nch W=10.8U L=0.34U
M27 PAD NVSS NVSS 0 nch W=24U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 GVSS TP4 Q 0 nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 GVSS TP13 TP4 0 nch W=4.1U L=0.24U
M33 TP20 TP0 VDD VDD pch W=3U L=0.24U
M34 TP20 TP0 GVSS 0 nch W=7U L=0.24U
R1I3234 N1I323TP7 EVSS 123
R1I3235 NVDD N1I323TP3 198
R1I3236 EVDD N1I323TP4 177
R1I3237 N1I323TP1 NVSS 198
R1I3238 N1I323TP5 NVSS 0.21
R1I3239 N1I323TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ciont25s3 DIN E PAD Q
C1I32810 PAD N1I328TP0 235FF
C1I32811 N1I328TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6U L=0.24U
M1I3280 N1I328TP7 N1I328TP0 NVDD NVDD pch W=38U L=0.34U
M1I3281 N1I328TP0 N1I328TP1 NVDD NVDD pch W=6U L=6U
M1I3282 N1I328TP2 N1I328TP3 NVSS NVSS nch W=6U L=6U
M1I3283 N1I328TP4 N1I328TP2 N1I328TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN GVSS 0 nch W=2U L=0.24U
M3 TP1 E VDD VDD pch W=6U L=0.24U
M4 TP1 E GVSS 0 nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=14U L=0.24U
M6 TP2 E TP3 0 nch W=10U L=0.24U
M7 TP3 TP1 GVSS 0 nch W=7.6U L=0.24U
M8 VDD TP20 TP2 VDD pch W=14U L=0.24U
M9 TP2 TP1 TP3 VDD pch W=10U L=0.24U
M10 GVSS TP20 TP3 0 nch W=7.6U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=84U L=0.34U
M14 TP14 TP3 NVSS 0 nch W=24.5U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=84U L=0.34U
M18 TP15 TP3 NVSS 0 nch W=24.5U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=84U L=0.34U
M22 TP16 TP3 NVSS 0 nch W=24.5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=84U L=0.34U
M26 TP17 TP3 NVSS 0 nch W=24.5U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 GVSS TP4 Q 0 nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 GVSS TP13 TP4 0 nch W=4.1U L=0.24U
M33 TP20 TP0 VDD VDD pch W=3U L=0.24U
M34 TP20 TP0 GVSS 0 nch W=7U L=0.24U
R1I3284 N1I328TP7 EVSS 123
R1I3285 NVDD N1I328TP3 198
R1I3286 EVDD N1I328TP4 177
R1I3287 N1I328TP1 NVSS 198
R1I3288 N1I328TP5 NVSS 0.21
R1I3289 N1I328TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ciont25s4 DIN E PAD Q
C1I32410 PAD N1I324TP0 235FF
C1I32411 N1I324TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6U L=0.24U
M1I3240 N1I324TP7 N1I324TP0 NVDD NVDD pch W=38U L=0.34U
M1I3241 N1I324TP0 N1I324TP1 NVDD NVDD pch W=6U L=6U
M1I3242 N1I324TP2 N1I324TP3 NVSS NVSS nch W=6U L=6U
M1I3243 N1I324TP4 N1I324TP2 N1I324TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN GVSS 0 nch W=2U L=0.24U
M3 TP20 E VDD VDD pch W=6U L=0.24U
M4 TP20 E GVSS 0 nch W=3U L=0.24U
M5 TP2 E VDD VDD pch W=18U L=0.24U
M6 TP2 E TP3 0 nch W=10U L=0.24U
M7 TP3 TP20 GVSS 0 nch W=10U L=0.24U
M8 VDD TP1 TP2 VDD pch W=18U L=0.24U
M9 TP2 TP20 TP3 VDD pch W=10U L=0.24U
M10 GVSS TP1 TP3 0 nch W=10U L=0.24U
M11 TP5 TP2 NVDD VDD pch W=152U L=0.34U
M14 TP14 TP3 NVSS 0 nch W=40.8U L=0.34U
M15 TP7 TP2 NVDD VDD pch W=152U L=0.34U
M18 TP15 TP3 NVSS 0 nch W=40.8U L=0.34U
M19 TP9 TP2 NVDD VDD pch W=152U L=0.34U
M22 TP16 TP3 NVSS 0 nch W=40.5U L=0.34U
M23 TP11 TP2 NVDD VDD pch W=152U L=0.34U
M26 TP17 TP3 NVSS 0 nch W=40.8U L=0.34U
M28 VDD TP4 Q VDD pch W=15.8U L=0.24U
M29 GVSS TP4 Q 0 nch W=8.8U L=0.24U
M30 VDD TP13 TP4 VDD pch W=5U L=0.24U
M31 GVSS TP13 TP4 0 nch W=4.1U L=0.24U
M33 TP1 TP0 VDD VDD pch W=3U L=0.24U
M34 TP1 TP0 GVSS 0 nch W=7U L=0.24U
R1I3244 N1I324TP7 EVSS 123
R1I3245 NVDD N1I324TP3 198
R1I3246 EVDD N1I324TP4 177
R1I3247 N1I324TP1 NVSS 198
R1I3248 N1I324TP5 NVSS 0.21
R1I3249 N1I324TP5 NVSS 0.21
R12 TP5 PAD 17
R16 TP7 PAD 17
R20 TP9 PAD 17
R24 TP11 PAD 17
R32 TP13 PAD 200
R34 PAD TP14 17
R35 PAD TP15 17
R36 PAD TP16 17
R37 PAD TP17 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_coi25s1 DIN PAD
C1I46610 PAD N1I466TP0 235FF
C1I46611 N1I466TP2 PAD 235FF
M1I4660 N1I466TP7 N1I466TP0 NVDD NVDD pch W=38U L=0.34U
M1I4661 N1I466TP0 N1I466TP1 NVDD NVDD pch W=6U L=6U
M1I4662 N1I466TP2 N1I466TP3 NVSS NVSS nch W=6U L=6U
M1I4663 N1I466TP4 N1I466TP2 N1I466TP5 NVSS nch W=38U L=0.34U
M3 TP1 DIN VDD VDD pch W=7.3U L=0.24U
M4 TP1 DIN GVSS 0 nch W=5.2U L=0.24U
M5 TP2 TP1 VDD VDD pch W=23.3U L=0.24U
M6 TP2 TP1 GVSS 0 nch W=9.2U L=0.24U
M7 TP3 TP2 NVDD VDD pch W=19U L=0.34U
M8 TP7 TP2 NVSS 0 nch W=6.5U L=0.34U
M9 TP4 TP2 NVDD VDD pch W=19U L=0.34U
M10 TP8 TP2 NVSS 0 nch W=6.5U L=0.34U
M11 TP5 TP2 NVDD VDD pch W=19U L=0.34U
M12 TP9 TP2 NVSS 0 nch W=6.5U L=0.34U
M13 TP6 TP2 NVDD VDD pch W=19U L=0.34U
M14 TP10 TP2 NVSS 0 nch W=6.5U L=0.34U
M15 PAD NVSS NVSS 0 nch W=20U L=0.34U
R1I4664 N1I466TP7 EVSS 123
R1I4665 NVDD N1I466TP3 198
R1I4666 EVDD N1I466TP4 177
R1I4667 N1I466TP1 NVSS 198
R1I4668 N1I466TP5 NVSS 0.21
R1I4669 N1I466TP5 NVSS 0.21
R15 TP3 PAD 17
R16 TP4 PAD 17
R17 TP5 PAD 17
R18 TP6 PAD 17
R19 PAD TP7 17
R20 PAD TP8 17
R21 PAD TP9 17
R22 PAD TP10 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_coi25s4 DIN PAD
C1I44310 PAD N1I443TP0 235FF
C1I44311 N1I443TP2 PAD 235FF
M1I4430 N1I443TP7 N1I443TP0 NVDD NVDD pch W=38U L=0.34U
M1I4431 N1I443TP0 N1I443TP1 NVDD NVDD pch W=6U L=6U
M1I4432 N1I443TP2 N1I443TP3 NVSS NVSS nch W=6U L=6U
M1I4433 N1I443TP4 N1I443TP2 N1I443TP5 NVSS nch W=38U L=0.34U
M3 TP1 DIN VDD VDD pch W=9.3U L=0.24U
M4 TP1 DIN GVSS 0 nch W=6.4U L=0.24U
M5 TP2 TP1 VDD VDD pch W=42.1U L=0.24U
M6 TP2 TP1 GVSS 0 nch W=17.2U L=0.24U
M7 TP3 TP2 NVDD VDD pch W=124U L=0.34U
M8 TP34 TP2 NVSS 0 nch W=40.5U L=0.34U
M9 TP31 TP2 NVDD VDD pch W=124U L=0.34U
M10 TP35 TP2 NVSS 0 nch W=40.5U L=0.34U
M11 TP32 TP2 NVDD VDD pch W=124U L=0.34U
M12 TP36 TP2 NVSS 0 nch W=40.5U L=0.34U
M13 TP33 TP2 NVDD VDD pch W=124U L=0.34U
M14 TP37 TP2 NVSS 0 nch W=40.5U L=0.34U
R1I4434 N1I443TP7 EVSS 123
R1I4435 NVDD N1I443TP3 198
R1I4436 EVDD N1I443TP4 177
R1I4437 N1I443TP1 NVSS 198
R1I4438 N1I443TP5 NVSS 0.21
R1I4439 N1I443TP5 NVSS 0.21
R15 TP3 PAD 17
R16 TP31 PAD 17
R17 TP32 PAD 17
R18 TP33 PAD 17
R19 PAD TP34 17
R20 PAD TP35 17
R21 PAD TP36 17
R22 PAD TP37 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_con25s1 DIN PAD
C1I46710 PAD N1I467TP0 235FF
C1I46711 N1I467TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6.2U L=0.24U
M1I4670 N1I467TP7 N1I467TP0 NVDD NVDD pch W=38U L=0.34U
M1I4671 N1I467TP0 N1I467TP1 NVDD NVDD pch W=6U L=6U
M1I4672 N1I467TP2 N1I467TP3 NVSS NVSS nch W=6U L=6U
M1I4673 N1I467TP4 N1I467TP2 N1I467TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN GVSS 0 nch W=3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=7.3U L=0.24U
M4 TP1 TP0 GVSS 0 nch W=5.2U L=0.24U
M5 TP2 TP1 VDD VDD pch W=23.3U L=0.24U
M6 TP2 TP1 GVSS 0 nch W=9.2U L=0.24U
M7 TP3 TP2 NVDD VDD pch W=19U L=0.34U
M8 TP7 TP2 NVSS 0 nch W=6.5U L=0.34U
M9 TP4 TP2 NVDD VDD pch W=19U L=0.34U
M10 TP8 TP2 NVSS 0 nch W=6.5U L=0.34U
M11 TP5 TP2 NVDD VDD pch W=19U L=0.34U
M12 TP9 TP2 NVSS 0 nch W=6.5U L=0.34U
M13 TP6 TP2 NVDD VDD pch W=19U L=0.34U
M14 TP10 TP2 NVSS 0 nch W=6.5U L=0.34U
M15 PAD NVSS NVSS 0 nch W=20U L=0.34U
R1I4674 N1I467TP7 EVSS 123
R1I4675 NVDD N1I467TP3 198
R1I4676 EVDD N1I467TP4 177
R1I4677 N1I467TP1 NVSS 198
R1I4678 N1I467TP5 NVSS 0.21
R1I4679 N1I467TP5 NVSS 0.21
R15 TP3 PAD 17
R16 TP4 PAD 17
R17 TP5 PAD 17
R18 TP6 PAD 17
R19 PAD TP7 17
R20 PAD TP8 17
R21 PAD TP9 17
R22 PAD TP10 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_con25s4 DIN PAD
C1I44410 PAD N1I444TP0 235FF
C1I44411 N1I444TP2 PAD 235FF
M1 TP0 DIN VDD VDD pch W=6.2U L=0.24U
M1I4440 N1I444TP7 N1I444TP0 NVDD NVDD pch W=38U L=0.34U
M1I4441 N1I444TP0 N1I444TP1 NVDD NVDD pch W=6U L=6U
M1I4442 N1I444TP2 N1I444TP3 NVSS NVSS nch W=6U L=6U
M1I4443 N1I444TP4 N1I444TP2 N1I444TP5 NVSS nch W=38U L=0.34U
M2 TP0 DIN GVSS 0 nch W=3U L=0.24U
M3 TP1 TP0 VDD VDD pch W=9.3U L=0.24U
M4 TP1 TP0 GVSS 0 nch W=6.4U L=0.24U
M5 TP2 TP1 VDD VDD pch W=42.1U L=0.24U
M6 TP2 TP1 GVSS 0 nch W=17.2U L=0.24U
M7 TP3 TP2 NVDD VDD pch W=124U L=0.34U
M8 TP34 TP2 NVSS 0 nch W=40.5U L=0.34U
M9 TP31 TP2 NVDD VDD pch W=124U L=0.34U
M10 TP35 TP2 NVSS 0 nch W=40.5U L=0.34U
M11 TP32 TP2 NVDD VDD pch W=124U L=0.34U
M12 TP36 TP2 NVSS 0 nch W=40.5U L=0.34U
M13 TP33 TP2 NVDD VDD pch W=124U L=0.34U
M14 TP37 TP2 NVSS 0 nch W=40.5U L=0.34U
R1I4444 N1I444TP7 EVSS 123
R1I4445 NVDD N1I444TP3 198
R1I4446 EVDD N1I444TP4 177
R1I4447 N1I444TP1 NVSS 198
R1I4448 N1I444TP5 NVSS 0.21
R1I4449 N1I444TP5 NVSS 0.21
R15 TP3 PAD 17
R16 TP31 PAD 17
R17 TP32 PAD 17
R18 TP33 PAD 17
R19 PAD TP34 17
R20 PAD TP35 17
R21 PAD TP36 17
R22 PAD TP37 17
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_corner INOUT2 INOUT1 AVCC AVSS VCC GVSS NVCC NVSS
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ncdavdd NVDD VDD AVDD EVDD PAD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 EVDD N1N43 NVSS NVSS nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N43 NVSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 NVDD PAD 0.0003
R3 AVDD VDD 0.0016
R4 VDD NVDD 0.0016
R5 EVDD PAD 0.0016
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ncdavss NVSS GVSS AVSS EVSS PAD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 EVSS N1N85 NVDD NVDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 NVDD N1N85 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 EVSS PAD 0.0024
R3 NVSS PAD 0.000966
R4 AVSS GVSS 0.002
R5 GVSS EVSS 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ncdvdd NVDD PAD VDD EVDD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 EVDD N1N43 NVSS NVSS nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N43 NVSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 NVDD PAD 0.003
R3 NVDD VDD 0.0016
R4 PAD EVDD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ncdvss NVSS PAD GVSS EVSS
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 GVSS N1N85 NVDD NVDD pch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 NVDD N1N85 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 EVSS PAD 0.002
R3 NVSS PAD 0.002
R4 GVSS EVSS 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ndavdd NVDD PAD AVDD EVDD
C1I2910 PAD N1I29TP0 235FF
C1I2911 N1I29TP2 PAD 235FF
M1 EVDD N1N44 NVSS NVSS nch W=300U L=0.34U
M1I290 N1I29TP7 N1I29TP0 NVDD NVDD pch W=38U L=0.34U
M1I291 N1I29TP0 N1I29TP1 NVDD NVDD pch W=6U L=6U
M1I292 N1I29TP2 N1I29TP3 NVSS NVSS nch W=6U L=6U
M1I293 N1I29TP4 N1I29TP2 N1I29TP5 NVSS nch W=38U L=0.34U
R1 N1N44 NVSS 400
R1I294 N1I29TP7 EVSS 123
R1I295 NVDD N1I29TP3 198
R1I296 EVDD N1I29TP4 177
R1I297 N1I29TP1 NVSS 198
R1I298 N1I29TP5 NVSS 0.21
R1I299 N1I29TP5 NVSS 0.21
R2 NVDD PAD 0.002
R3 AVDD NVDD 0.002
R4 EVDD PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ndavss NVSS PAD EVSS AVSS
C1I6210 PAD N1I62TP0 235FF
C1I6211 N1I62TP2 PAD 235FF
M1 EVSS N1N56 NVDD NVDD pch W=300U L=0.34U
M1I620 N1I62TP7 N1I62TP0 NVDD NVDD pch W=38U L=0.34U
M1I621 N1I62TP0 N1I62TP1 NVDD NVDD pch W=6U L=6U
M1I622 N1I62TP2 N1I62TP3 NVSS NVSS nch W=6U L=6U
M1I623 N1I62TP4 N1I62TP2 N1I62TP5 NVSS nch W=38U L=0.34U
R1 NVDD N1N56 400
R1I624 N1I62TP7 EVSS 123
R1I625 NVDD N1I62TP3 198
R1I626 EVDD N1I62TP4 177
R1I627 N1I62TP1 NVSS 198
R1I628 N1I62TP5 NVSS 0.21
R1I629 N1I62TP5 NVSS 0.21
R2 EVSS PAD 0.001
R3 NVSS PAD 0.00035
R4 AVSS EVSS 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ndvdd EVDD NVDD PAD N1
C1I6210 PAD N1I62TP0 235FF
C1I6211 N1I62TP2 PAD 235FF
M1 EVDD N1N44 NVSS NVSS nch W=300U L=0.34U
M1I620 N1I62TP7 N1I62TP0 NVDD NVDD pch W=38U L=0.34U
M1I621 N1I62TP0 N1I62TP1 NVDD NVDD pch W=6U L=6U
M1I622 N1I62TP2 N1I62TP3 NVSS NVSS nch W=6U L=6U
M1I623 N1I62TP4 N1I62TP2 N1I62TP5 NVSS nch W=38U L=0.34U
R1 N1N44 NVSS 400
R1I624 N1I62TP7 EVSS 123
R1I625 NVDD N1I62TP3 198
R1I626 EVDD N1I62TP4 177
R1I627 N1I62TP1 NVSS 198
R1I628 N1I62TP5 NVSS 0.21
R1I629 N1I62TP5 NVSS 0.21
R2 NVDD PAD 0.0023
R3 PAD EVDD 0.0018
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT gated_ndvss NVSS PAD EVSS N1
C1I6210 PAD N1I62TP0 235FF
C1I6211 N1I62TP2 PAD 235FF
M1 EVSS N1N56 NVDD NVDD pch W=300U L=0.34U
M1I620 N1I62TP7 N1I62TP0 NVDD NVDD pch W=38U L=0.34U
M1I621 N1I62TP0 N1I62TP1 NVDD NVDD pch W=6U L=6U
M1I622 N1I62TP2 N1I62TP3 NVSS NVSS nch W=6U L=6U
M1I623 N1I62TP4 N1I62TP2 N1I62TP5 NVSS nch W=38U L=0.34U
R1 NVDD N1N56 400
R1I624 N1I62TP7 EVSS 123
R1I625 NVDD N1I62TP3 198
R1I626 EVDD N1I62TP4 177
R1I627 N1I62TP1 NVSS 198
R1I628 N1I62TP5 NVSS 0.21
R1I629 N1I62TP5 NVSS 0.21
R2 NVSS PAD 0.0027
R3 EVSS PAD 0.002
.GLOBAL VDD
.GLOBAL VSS
.ENDS

.SUBCKT and9s1 DIN1 DIN2 DIN3 DIN4 DIN5 DIN6 DIN7 DIN8 DIN9 Q
M5 N1N304 DIN1 N1N314 VSS nch W=6.3U L=0.24U
M1 N1N304 DIN1 VDD VDD pch W=2.1U L=0.24U
M2 N1N304 DIN2 VDD VDD pch W=2.1U L=0.24U
M3 N1N304 DIN3 VDD VDD pch W=2.1U L=0.24U
M4 N1N304 DIN4 VDD VDD pch W=2.1U L=0.24U
M6 N1N314 DIN2 N1N316 VSS nch W=6.5U L=0.24U
M7 N1N316 DIN3 N1N318 VSS nch W=6.7U L=0.24U
M8 N1N318 DIN4 VSS VSS nch W=6.9U L=0.24U
M9 N1N343 N1N304 VDD VDD pch W=5.4U L=0.24U
M10 N1N343 N1N413 N1N345 VDD pch W=5.4U L=0.24U
M11 N1N345 N1N304 VSS VSS nch W=1.5U L=0.24U
M12 VSS N1N413 N1N345 VSS nch W=1.5U L=0.24U
M13 N1N413 DIN5 VDD VDD pch W=2.1U L=0.24U
M14 N1N413 DIN6 VDD VDD pch W=2.1U L=0.24U
M15 N1N413 DIN7 VDD VDD pch W=2.1U L=0.24U
M16 N1N413 DIN8 VDD VDD pch W=2.1U L=0.24U
M17 N1N413 DIN5 N1N362 VSS nch W=6.3U L=0.24U
M18 N1N362 DIN6 N1N364 VSS nch W=6.5U L=0.24U
M19 N1N364 DIN7 N1N366 VSS nch W=6.7U L=0.24U
M20 N1N366 DIN8 VSS VSS nch W=6.9U L=0.24U
M22 Q N1N345 VSS VSS nch W=3U L=0.24U
M21 Q N1N345 VDD VDD pch W=6.5U L=0.24U
.GLOBAL VDD
.GLOBAL VSS
.ENDS
