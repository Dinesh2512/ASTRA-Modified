module sha256(
    input [511:0] block,
    input clk,
    input rst,
    input init,
    input next,
    input sel,
    output [255:0] digest,
    output ready,
    output digest_valid,
    output [15:0] pufout);

    wire n1755, n1747, n1754, n1752, n1751, n1750, n1749, n1748, n1753, n1746, n1745, n1651, n1650, n1682, n1649, n1681, n1648, n1680, n1647, n1679;
    wire n1646, n1678, n1645, n1677, n1644, n1676, n1643, n1675, n1642, n1674, n1641, n1673, n1640, n1672, n1639, n1671, n1638, n1670, n1637, n1669;
    wire n1636, n1668, n1635, n1667, n1634, n1666, n1633, n1665, n1632, n1664, n1631, n1663, n1630, n1662, n1629, n1661, n1628, n1660, n1627, n1659;
    wire n1626, n1658, n1625, n1657, n1624, n1656, n1623, n1655, n1622, n1654, n1621, n1653, n1620, n1652, n1619, n1587, n1586, n1618, n1585, n1617;
    wire n1584, n1616, n1583, n1615, n1582, n1614, n1581, n1613, n1580, n1612, n1579, n1611, n1578, n1610, n1577, n1609, n1576, n1608, n1575, n1607;
    wire n1574, n1606, n1573, n1605, n1572, n1604, n1571, n1603, n1570, n1602, n1569, n1601, n1568, n1600, n1567, n1599, n1566, n1598, n1565, n1597;
    wire n1564, n1596, n1563, n1595, n1562, n1594, n1561, n1593, n1560, n1592, n1559, n1591, n1558, n1590, n1557, n1589, n1556, n1588, n1555, n1523;
    wire n1522, n1554, n1521, n1553, n1520, n1552, n1519, n1551, n1518, n1550, n1517, n1549, n1516, n1548, n1515, n1547, n1514, n1546, n1513, n1545;
    wire n1512, n1544, n1511, n1543, n1510, n1542, n1509, n1541, n1508, n1540, n1507, n1539, n1506, n1538, n1505, n1537, n1504, n1536, n1503, n1535;
    wire n1502, n1534, n1501, n1533, n1500, n1532, n1499, n1531, n1498, n1530, n1497, n1529, n1496, n1528, n1495, n1527, n1494, n1526, n1493, n1525;
    wire n1492, n1524, n1491, n1459, n1458, n1490, n1457, n1489, n1456, n1488, n1455, n1487, n1454, n1486, n1453, n1485, n1452, n1484, n1451, n1483;
    wire n1450, n1482, n1449, n1481, n1448, n1480, n1447, n1479, n1446, n1478, n1445, n1477, n1444, n1476, n1443, n1475, n1442, n1474, n1441, n1473;
    wire n1440, n1472, n1439, n1471, n1438, n1470, n1437, n1469, n1436, n1468, n1435, n1467, n1434, n1466, n1433, n1465, n1432, n1464, n1431, n1463;
    wire n1430, n1462, n1429, n1461, n1428, n1460, n1427, n1395, n1394, n1426, n1393, n1425, n1392, n1424, n1391, n1423, n1390, n1422, n1389, n1421;
    wire n1388, n1420, n1387, n1419, n1386, n1418, n1385, n1417, n1384, n1416, n1383, n1415, n1382, n1414, n1381, n1413, n1380, n1412, n1379, n1411;
    wire n1378, n1410, n1377, n1409, n1376, n1408, n1375, n1407, n1374, n1406, n1373, n1405, n1372, n1404, n1371, n1403, n1370, n1402, n1369, n1401;
    wire n1368, n1400, n1367, n1399, n1366, n1398, n1365, n1397, n1364, n1396, n1363, n1331, n1330, n1362, n1329, n1361, n1328, n1360, n1327, n1359;
    wire n1326, n1358, n1325, n1357, n1324, n1356, n1323, n1355, n1322, n1354, n1321, n1353, n1320, n1352, n1319, n1351, n1318, n1350, n1317, n1349;
    wire n1316, n1348, n1315, n1347, n1314, n1346, n1313, n1345, n1312, n1344, n1311, n1343, n1310, n1342, n1309, n1341, n1308, n1340, n1307, n1339;
    wire n1306, n1338, n1305, n1337, n1304, n1336, n1303, n1335, n1302, n1334, n1301, n1333, n1300, n1332, n1299, n1267, n1266, n1298, n1265, n1297;
    wire n1264, n1296, n1263, n1295, n1262, n1294, n1261, n1293, n1260, n1292, n1259, n1291, n1258, n1290, n1257, n1289, n1256, n1288, n1255, n1287;
    wire n1254, n1286, n1253, n1285, n1252, n1284, n1251, n1283, n1250, n1282, n1249, n1281, n1248, n1280, n1247, n1279, n1246, n1278, n1245, n1277;
    wire n1244, n1276, n1243, n1275, n1242, n1274, n1241, n1273, n1240, n1272, n1239, n1271, n1238, n1270, n1237, n1269, n1236, n1268, n1235, n1714;
    wire n1713, n1744, n1712, n1743, n1711, n1742, n1710, n1741, n1709, n1740, n1708, n1739, n1707, n1738, n1706, n1737, n1705, n1736, n1704, n1735;
    wire n1703, n1734, n1702, n1733, n1701, n1732, n1700, n1731, n1699, n1730, n1698, n1729, n1697, n1728, n1696, n1727, n1695, n1726, n1694, n1725;
    wire n1693, n1724, n1692, n1723, n1691, n1722, n1690, n1721, n1689, n1720, n1688, n1719, n1687, n1718, n1686, n1717, n1685, n1716, n1684, n1715;
    wire n1683, w_mem_inst_n1624, w_mem_inst_n1656, w_mem_inst_n1688, w_mem_inst_n1720, w_mem_inst_n1752, w_mem_inst_n1784, w_mem_inst_n1816, w_mem_inst_n1848, w_mem_inst_n1880, w_mem_inst_n1912, w_mem_inst_n1944, w_mem_inst_n1976, w_mem_inst_n2008, w_mem_inst_n2040, w_mem_inst_n2072, w_mem_inst_n2104, w_mem_inst_n1625, w_mem_inst_n1657, w_mem_inst_n1689;
    wire w_mem_inst_n1721, w_mem_inst_n1753, w_mem_inst_n1785, w_mem_inst_n1817, w_mem_inst_n1849, w_mem_inst_n1881, w_mem_inst_n1913, w_mem_inst_n1945, w_mem_inst_n1977, w_mem_inst_n2009, w_mem_inst_n2041, w_mem_inst_n2073, w_mem_inst_n2105, w_mem_inst_n1626, w_mem_inst_n1658, w_mem_inst_n1690, w_mem_inst_n1722, w_mem_inst_n1754, w_mem_inst_n1786, w_mem_inst_n1818;
    wire w_mem_inst_n1850, w_mem_inst_n1882, w_mem_inst_n1914, w_mem_inst_n1946, w_mem_inst_n1978, w_mem_inst_n2010, w_mem_inst_n2042, w_mem_inst_n2074, w_mem_inst_n2106, w_mem_inst_n1627, w_mem_inst_n1659, w_mem_inst_n1691, w_mem_inst_n1723, w_mem_inst_n1755, w_mem_inst_n1787, w_mem_inst_n1819, w_mem_inst_n1851, w_mem_inst_n1883, w_mem_inst_n1915, w_mem_inst_n1947;
    wire w_mem_inst_n1979, w_mem_inst_n2011, w_mem_inst_n2043, w_mem_inst_n2075, w_mem_inst_n2107, w_mem_inst_n1628, w_mem_inst_n1660, w_mem_inst_n1692, w_mem_inst_n1724, w_mem_inst_n1756, w_mem_inst_n1788, w_mem_inst_n1820, w_mem_inst_n1852, w_mem_inst_n1884, w_mem_inst_n1916, w_mem_inst_n1948, w_mem_inst_n1980, w_mem_inst_n2012, w_mem_inst_n2044, w_mem_inst_n2076;
    wire w_mem_inst_n2108, w_mem_inst_n1629, w_mem_inst_n1661, w_mem_inst_n1693, w_mem_inst_n1725, w_mem_inst_n1757, w_mem_inst_n1789, w_mem_inst_n1821, w_mem_inst_n1853, w_mem_inst_n1885, w_mem_inst_n1917, w_mem_inst_n1949, w_mem_inst_n1981, w_mem_inst_n2013, w_mem_inst_n2045, w_mem_inst_n2077, w_mem_inst_n2109, w_mem_inst_n1630, w_mem_inst_n1662, w_mem_inst_n1694;
    wire w_mem_inst_n1726, w_mem_inst_n1758, w_mem_inst_n1790, w_mem_inst_n1822, w_mem_inst_n1854, w_mem_inst_n1886, w_mem_inst_n1918, w_mem_inst_n1950, w_mem_inst_n1982, w_mem_inst_n2014, w_mem_inst_n2046, w_mem_inst_n2078, w_mem_inst_n2110, w_mem_inst_n1631, w_mem_inst_n1663, w_mem_inst_n1695, w_mem_inst_n1727, w_mem_inst_n1759, w_mem_inst_n1791, w_mem_inst_n1823;
    wire w_mem_inst_n1855, w_mem_inst_n1887, w_mem_inst_n1919, w_mem_inst_n1951, w_mem_inst_n1983, w_mem_inst_n2015, w_mem_inst_n2047, w_mem_inst_n2079, w_mem_inst_n2111, w_mem_inst_n1632, w_mem_inst_n1664, w_mem_inst_n1696, w_mem_inst_n1728, w_mem_inst_n1760, w_mem_inst_n1792, w_mem_inst_n1824, w_mem_inst_n1856, w_mem_inst_n1888, w_mem_inst_n1920, w_mem_inst_n1952;
    wire w_mem_inst_n1984, w_mem_inst_n2016, w_mem_inst_n2048, w_mem_inst_n2080, w_mem_inst_n2112, w_mem_inst_n1633, w_mem_inst_n1665, w_mem_inst_n1697, w_mem_inst_n1729, w_mem_inst_n1761, w_mem_inst_n1793, w_mem_inst_n1825, w_mem_inst_n1857, w_mem_inst_n1889, w_mem_inst_n1921, w_mem_inst_n1953, w_mem_inst_n1985, w_mem_inst_n2017, w_mem_inst_n2049, w_mem_inst_n2081;
    wire w_mem_inst_n2113, w_mem_inst_n1634, w_mem_inst_n1666, w_mem_inst_n1698, w_mem_inst_n1730, w_mem_inst_n1762, w_mem_inst_n1794, w_mem_inst_n1826, w_mem_inst_n1858, w_mem_inst_n1890, w_mem_inst_n1922, w_mem_inst_n1954, w_mem_inst_n1986, w_mem_inst_n2018, w_mem_inst_n2050, w_mem_inst_n2082, w_mem_inst_n2114, w_mem_inst_n1635, w_mem_inst_n1667, w_mem_inst_n1699;
    wire w_mem_inst_n1731, w_mem_inst_n1763, w_mem_inst_n1795, w_mem_inst_n1827, w_mem_inst_n1859, w_mem_inst_n1891, w_mem_inst_n1923, w_mem_inst_n1955, w_mem_inst_n1987, w_mem_inst_n2019, w_mem_inst_n2051, w_mem_inst_n2083, w_mem_inst_n2115, w_mem_inst_n1636, w_mem_inst_n1668, w_mem_inst_n1700, w_mem_inst_n1732, w_mem_inst_n1764, w_mem_inst_n1796, w_mem_inst_n1828;
    wire w_mem_inst_n1860, w_mem_inst_n1892, w_mem_inst_n1924, w_mem_inst_n1956, w_mem_inst_n1988, w_mem_inst_n2020, w_mem_inst_n2052, w_mem_inst_n2084, w_mem_inst_n2116, w_mem_inst_n1637, w_mem_inst_n1669, w_mem_inst_n1701, w_mem_inst_n1733, w_mem_inst_n1765, w_mem_inst_n1797, w_mem_inst_n1829, w_mem_inst_n1861, w_mem_inst_n1893, w_mem_inst_n1925, w_mem_inst_n1957;
    wire w_mem_inst_n1989, w_mem_inst_n2021, w_mem_inst_n2053, w_mem_inst_n2085, w_mem_inst_n2117, w_mem_inst_n1638, w_mem_inst_n1670, w_mem_inst_n1702, w_mem_inst_n1734, w_mem_inst_n1766, w_mem_inst_n1798, w_mem_inst_n1830, w_mem_inst_n1862, w_mem_inst_n1894, w_mem_inst_n1926, w_mem_inst_n1958, w_mem_inst_n1990, w_mem_inst_n2022, w_mem_inst_n2054, w_mem_inst_n2086;
    wire w_mem_inst_n2118, w_mem_inst_n1639, w_mem_inst_n1671, w_mem_inst_n1703, w_mem_inst_n1735, w_mem_inst_n1767, w_mem_inst_n1799, w_mem_inst_n1831, w_mem_inst_n1863, w_mem_inst_n1895, w_mem_inst_n1927, w_mem_inst_n1959, w_mem_inst_n1991, w_mem_inst_n2023, w_mem_inst_n2055, w_mem_inst_n2087, w_mem_inst_n2119, w_mem_inst_n1640, w_mem_inst_n1672, w_mem_inst_n1704;
    wire w_mem_inst_n1736, w_mem_inst_n1768, w_mem_inst_n1800, w_mem_inst_n1832, w_mem_inst_n1864, w_mem_inst_n1896, w_mem_inst_n1928, w_mem_inst_n1960, w_mem_inst_n1992, w_mem_inst_n2024, w_mem_inst_n2056, w_mem_inst_n2088, w_mem_inst_n2120, w_mem_inst_n1641, w_mem_inst_n1673, w_mem_inst_n1705, w_mem_inst_n1737, w_mem_inst_n1769, w_mem_inst_n1801, w_mem_inst_n1833;
    wire w_mem_inst_n1865, w_mem_inst_n1897, w_mem_inst_n1929, w_mem_inst_n1961, w_mem_inst_n1993, w_mem_inst_n2025, w_mem_inst_n2057, w_mem_inst_n2089, w_mem_inst_n2121, w_mem_inst_n1642, w_mem_inst_n1674, w_mem_inst_n1706, w_mem_inst_n1738, w_mem_inst_n1770, w_mem_inst_n1802, w_mem_inst_n1834, w_mem_inst_n1866, w_mem_inst_n1898, w_mem_inst_n1930, w_mem_inst_n1962;
    wire w_mem_inst_n1994, w_mem_inst_n2026, w_mem_inst_n2058, w_mem_inst_n2090, w_mem_inst_n2122, w_mem_inst_n1643, w_mem_inst_n1675, w_mem_inst_n1707, w_mem_inst_n1739, w_mem_inst_n1771, w_mem_inst_n1803, w_mem_inst_n1835, w_mem_inst_n1867, w_mem_inst_n1899, w_mem_inst_n1931, w_mem_inst_n1963, w_mem_inst_n1995, w_mem_inst_n2027, w_mem_inst_n2059, w_mem_inst_n2091;
    wire w_mem_inst_n2123, w_mem_inst_n1644, w_mem_inst_n1676, w_mem_inst_n1708, w_mem_inst_n1740, w_mem_inst_n1772, w_mem_inst_n1804, w_mem_inst_n1836, w_mem_inst_n1868, w_mem_inst_n1900, w_mem_inst_n1932, w_mem_inst_n1964, w_mem_inst_n1996, w_mem_inst_n2028, w_mem_inst_n2060, w_mem_inst_n2092, w_mem_inst_n2124, w_mem_inst_n1645, w_mem_inst_n1677, w_mem_inst_n1709;
    wire w_mem_inst_n1741, w_mem_inst_n1773, w_mem_inst_n1805, w_mem_inst_n1837, w_mem_inst_n1869, w_mem_inst_n1901, w_mem_inst_n1933, w_mem_inst_n1965, w_mem_inst_n1997, w_mem_inst_n2029, w_mem_inst_n2061, w_mem_inst_n2093, w_mem_inst_n2125, w_mem_inst_n1646, w_mem_inst_n1678, w_mem_inst_n1710, w_mem_inst_n1742, w_mem_inst_n1774, w_mem_inst_n1806, w_mem_inst_n1838;
    wire w_mem_inst_n1870, w_mem_inst_n1902, w_mem_inst_n1934, w_mem_inst_n1966, w_mem_inst_n1998, w_mem_inst_n2030, w_mem_inst_n2062, w_mem_inst_n2094, w_mem_inst_n2126, w_mem_inst_n1647, w_mem_inst_n1679, w_mem_inst_n1711, w_mem_inst_n1743, w_mem_inst_n1775, w_mem_inst_n1807, w_mem_inst_n1839, w_mem_inst_n1871, w_mem_inst_n1903, w_mem_inst_n1935, w_mem_inst_n1967;
    wire w_mem_inst_n1999, w_mem_inst_n2031, w_mem_inst_n2063, w_mem_inst_n2095, w_mem_inst_n2127, w_mem_inst_n1648, w_mem_inst_n1680, w_mem_inst_n1712, w_mem_inst_n1744, w_mem_inst_n1776, w_mem_inst_n1808, w_mem_inst_n1840, w_mem_inst_n1872, w_mem_inst_n1904, w_mem_inst_n1936, w_mem_inst_n1968, w_mem_inst_n2000, w_mem_inst_n2032, w_mem_inst_n2064, w_mem_inst_n2096;
    wire w_mem_inst_n2128, w_mem_inst_n1649, w_mem_inst_n1681, w_mem_inst_n1713, w_mem_inst_n1745, w_mem_inst_n1777, w_mem_inst_n1809, w_mem_inst_n1841, w_mem_inst_n1873, w_mem_inst_n1905, w_mem_inst_n1937, w_mem_inst_n1969, w_mem_inst_n2001, w_mem_inst_n2033, w_mem_inst_n2065, w_mem_inst_n2097, w_mem_inst_n2129, w_mem_inst_n1650, w_mem_inst_n1682, w_mem_inst_n1714;
    wire w_mem_inst_n1746, w_mem_inst_n1778, w_mem_inst_n1810, w_mem_inst_n1842, w_mem_inst_n1874, w_mem_inst_n1906, w_mem_inst_n1938, w_mem_inst_n1970, w_mem_inst_n2002, w_mem_inst_n2034, w_mem_inst_n2066, w_mem_inst_n2098, w_mem_inst_n2130, w_mem_inst_n1651, w_mem_inst_n1683, w_mem_inst_n1715, w_mem_inst_n1747, w_mem_inst_n1779, w_mem_inst_n1811, w_mem_inst_n1843;
    wire w_mem_inst_n1875, w_mem_inst_n1907, w_mem_inst_n1939, w_mem_inst_n1971, w_mem_inst_n2003, w_mem_inst_n2035, w_mem_inst_n2067, w_mem_inst_n2099, w_mem_inst_n2131, w_mem_inst_n1652, w_mem_inst_n1684, w_mem_inst_n1716, w_mem_inst_n1748, w_mem_inst_n1780, w_mem_inst_n1812, w_mem_inst_n1844, w_mem_inst_n1876, w_mem_inst_n1908, w_mem_inst_n1940, w_mem_inst_n1972;
    wire w_mem_inst_n2004, w_mem_inst_n2036, w_mem_inst_n2068, w_mem_inst_n2100, w_mem_inst_n2132, w_mem_inst_n1653, w_mem_inst_n1685, w_mem_inst_n1717, w_mem_inst_n1749, w_mem_inst_n1781, w_mem_inst_n1813, w_mem_inst_n1845, w_mem_inst_n1877, w_mem_inst_n1909, w_mem_inst_n1941, w_mem_inst_n1973, w_mem_inst_n2005, w_mem_inst_n2037, w_mem_inst_n2069, w_mem_inst_n2101;
    wire w_mem_inst_n2133, w_mem_inst_n1654, w_mem_inst_n1686, w_mem_inst_n1718, w_mem_inst_n1750, w_mem_inst_n1782, w_mem_inst_n1814, w_mem_inst_n1846, w_mem_inst_n1878, w_mem_inst_n1910, w_mem_inst_n1942, w_mem_inst_n1974, w_mem_inst_n2006, w_mem_inst_n2038, w_mem_inst_n2070, w_mem_inst_n2102, w_mem_inst_n2134, w_mem_inst_n1655, w_mem_inst_n1687, w_mem_inst_n1719;
    wire w_mem_inst_n1751, w_mem_inst_n1783, w_mem_inst_n1815, w_mem_inst_n1847, w_mem_inst_n1879, w_mem_inst_n1911, w_mem_inst_n1943, w_mem_inst_n1975, w_mem_inst_n2007, w_mem_inst_n2039, w_mem_inst_n2071, w_mem_inst_n2103, w_mem_inst_n2135, w_mem_inst_n2136, w_mem_inst_n2137, w_mem_inst_n2138, w_mem_inst_n2139, w_mem_inst_n2141, w_mem_inst_sha256_w_mem_ctrl_reg_0_, w_mem_inst_n2140;
    wire w_mem_inst_n2142, w_mem_inst_N641, w_mem_inst_N638, n2964, w_mem_inst_N642, w_mem_inst_N637, w_mem_inst_N643, w_mem_inst_N636, w_mem_inst_N644, w_mem_inst_N635, w_mem_inst_N645, w_mem_inst_N634, w_mem_inst_N646, w_mem_inst_N633, w_mem_inst_N647, w_mem_inst_N632, w_mem_inst_N648, w_mem_inst_N631, w_mem_inst_N649, w_mem_inst_N630;
    wire w_mem_inst_N650, w_mem_inst_N629, w_mem_inst_N651, w_mem_inst_N628, w_mem_inst_N652, w_mem_inst_N627, w_mem_inst_N653, w_mem_inst_N626, w_mem_inst_N654, w_mem_inst_N625, w_mem_inst_N655, w_mem_inst_N624, w_mem_inst_N656, w_mem_inst_N623, w_mem_inst_N657, w_mem_inst_N622, w_mem_inst_N658, w_mem_inst_N621, w_mem_inst_N659, w_mem_inst_N620;
    wire w_mem_inst_N660, w_mem_inst_N619, w_mem_inst_N661, w_mem_inst_N618, w_mem_inst_N662, w_mem_inst_N617, w_mem_inst_N663, w_mem_inst_N616, w_mem_inst_N664, w_mem_inst_N615, w_mem_inst_N665, w_mem_inst_N614, w_mem_inst_N666, w_mem_inst_N613, w_mem_inst_N667, w_mem_inst_N612, w_mem_inst_N668, w_mem_inst_N611, w_mem_inst_N669, w_mem_inst_N610;
    wire w_mem_inst_N670, w_mem_inst_N609, w_mem_inst_N671, w_mem_inst_N608, w_mem_inst_N673, w_mem_inst_N606, n2965, w_mem_inst_N674, w_mem_inst_N605, w_mem_inst_N675, w_mem_inst_N604, w_mem_inst_N676, w_mem_inst_N603, w_mem_inst_N677, w_mem_inst_N602, w_mem_inst_N678, w_mem_inst_N601, w_mem_inst_N679, w_mem_inst_N600, w_mem_inst_N680;
    wire w_mem_inst_N599, w_mem_inst_N681, w_mem_inst_N598, w_mem_inst_N682, w_mem_inst_N597, w_mem_inst_N683, w_mem_inst_N596, w_mem_inst_N684, w_mem_inst_N595, w_mem_inst_N685, w_mem_inst_N594, w_mem_inst_N686, w_mem_inst_N593, w_mem_inst_N687, w_mem_inst_N592, w_mem_inst_N688, w_mem_inst_N591, w_mem_inst_N689, w_mem_inst_N590, w_mem_inst_N690;
    wire w_mem_inst_N589, w_mem_inst_N691, w_mem_inst_N588, w_mem_inst_N692, w_mem_inst_N587, w_mem_inst_N693, w_mem_inst_N586, w_mem_inst_N694, w_mem_inst_N585, w_mem_inst_N695, w_mem_inst_N584, w_mem_inst_N696, w_mem_inst_N583, w_mem_inst_N697, w_mem_inst_N582, w_mem_inst_N698, w_mem_inst_N581, w_mem_inst_N699, w_mem_inst_N580, w_mem_inst_N700;
    wire w_mem_inst_N579, w_mem_inst_N701, w_mem_inst_N578, w_mem_inst_N702, w_mem_inst_N577, w_mem_inst_N703, w_mem_inst_N576, n2962, w_mem_inst_N711, w_mem_inst_N712, w_mem_inst_N713, w_mem_inst_N714, N1615, N1616, N1617, N1618, N1580, n2967, N1581, N1582;
    wire N1583, N1584, N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594, N1595, N1596, N1597, N1598, N1599, N1600, N1601, N1602;
    wire N1603, N1604, N1605, N1606, N1607, N1608, N1609, N1610, N1548, N1028, n2960, N1549, n6194, N1550, N1026, N1551, N1025, N1552, N1024, N1553;
    wire N1023, N1554, N1022, N1555, N1021, N1556, n6195, N1557, n6196, N1558, N1018, N1559, N1017, N1560, N1016, N1561, N1015, N1562, N1014, N1563;
    wire N1013, N1564, N1012, N1565, N1011, N1566, N1010, N1567, N1009, N1568, N1008, N1569, N1007, N1570, N1006, N1571, N1005, N1572, n6197, N1573;
    wire N1003, N1574, n6198, N1575, N1001, N1576, n6199, N1577, N999, N1578, N998, N996, n2963, N995, N994, N993, N992, N991, N990, N989;
    wire N988, N987, N986, N985, N984, N983, N982, N981, N980, N979, N978, N977, N976, N975, N974, N973, N972, N971, N970, N969;
    wire N968, N967, N966, N903, N935, n2959, N904, N936, N905, N937, N906, N938, N907, N939, N908, N940, N909, N941, N910, N942;
    wire N911, N943, N912, N944, N913, N945, N914, N946, N915, N947, N916, N948, N917, N949, N918, N950, N919, N951, N920, N952;
    wire N921, N953, N922, N954, N923, N955, N924, N956, N925, N957, N926, N958, N927, N959, N928, N960, N929, N961, N930, N962;
    wire N931, N963, N932, N964, N933, N965, n1818, N871, n2961, n1774, N872, n1773, N873, n1772, N874, n1771, N875, N876, N877, n1770;
    wire N878, n1769, N879, n1768, N880, n2779, N881, N882, n1767, N883, n1817, N884, n2086, N885, n1766, N886, N887, n1765, N888, N889;
    wire n2649, N890, n1764, N891, n1763, N892, n2072, N893, n1762, N894, n2537, N895, n2480, N896, n1761, N897, n1760, N898, N899, N900;
    wire n1816, N901, N868, n1757, n1850, N867, n1848, N866, n1847, N865, n1846, N864, n1845, N863, n1844, N862, n1843, N861, n1842, N860;
    wire n1841, N859, n1830, N858, n1829, N857, n1828, N856, n1827, N855, n1826, N854, n1825, N853, n1824, N852, n1823, N851, n1822, N850;
    wire n1821, N849, n1820, N848, n1819, N847, n1840, N846, n1839, N845, n1838, N844, n1837, N843, n1836, N842, n1835, N841, n1834, N840;
    wire n1833, N839, n1832, N838, n1831, N836, n2966, N835, N834, N833, N832, N831, N830, N829, N828, N827, N826, N825, N824, N823;
    wire N822, N821, N820, N819, N818, N817, N816, N815, N814, N813, N812, N811, N810, N809, N808, N807, N806, N775, n2969, N776;
    wire N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796;
    wire N797, N798, N799, N800, N801, N802, N803, N804, N805, N743, n2974, N744, N745, N746, N747, N748, N749, N750, N751, N752;
    wire N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772;
    wire N773, N711, n2970, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726, N727, N728;
    wire N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N679, n2975, N680, N681, N682, N683, N684;
    wire N685, N686, N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704;
    wire N705, N706, N707, N708, N709, N647, n2971, N648, N649, N650, N651, N652, N653, N654, N655, N656, N657, N658, N659, N660;
    wire N661, N662, N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N615, n2972, N616;
    wire N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636;
    wire N637, N638, N639, N640, N641, N642, N643, N644, N645, N583, n2968, N584, N585, N586, N587, N588, N589, N590, N591, N592;
    wire N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612;
    wire N613, N551, n2973, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568;
    wire N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, n5971, n2718, n2595, n5991, n5821, n2893, n5770;
    wire n2847, n2783, n5751, n2657, n2720, n5749, n2890, n2107, n6033, n2845, n5837, n5839, n2712, n4169, n2894, n2958, n5853, n2955, n2717, n4170;
    wire n4442, n1953, n5752, n5771, n5793, n5786, n5867, n5843, n3103, n2777, n3100, n1756, n5912, n1777, n2023, n1778, n1758, n2100, n1776, n4783;
    wire n2951, n4713, n1759, n2127, n1780, n2065, n1866, n2068, n1867, n2071, n1858, n2074, n1856, n2077, n1859, n2082, n1860, n2085, n1865, n2091;
    wire n1868, n2094, n1869, n2046, n1861, n2048, n1855, n2051, n1862, n2054, n1863, n2057, n1864, n2062, n1857, n5848, n2891, n5861, n2849, n1775;
    wire n1936, n1854, n2099, n1871, n1877, n5981, n1898, n2022, n1779, n1941, n1875, n3115, n1781, n1974, n1872, n1782, n1878, n1982, n1783, n1879;
    wire n1984, n1784, n1880, n1986, n1785, n1881, n1988, n1786, n1882, n1990, n1787, n1883, n1992, n1788, n1884, n1994, n1789, n1885, n1996, n1790;
    wire n1886, n1998, n1791, n1887, n2000, n1792, n1888, n2002, n1793, n1889, n2004, n1794, n1890, n2006, n1795, n1891, n2008, n1796, n1892, n2010;
    wire n1797, n1893, n2012, n1798, n1894, n2014, n1799, n1895, n2016, n1800, n1896, n2018, n1801, n1897, n2020, n1802, n1899, n2024, n1803, n1900;
    wire n2026, n1804, n1901, n2028, n1805, n1902, n2030, n1806, n1903, n2032, n1807, n1904, n2034, n1808, n1905, n2036, n1809, n1906, n2038, n1810;
    wire n1907, n2040, n1811, n1908, n2042, n1812, n1876, n2095, n1813, n1874, n2078, n1814, n1873, n2087, n1815, n2058, n1870, n2059, n2088, n2079;
    wire n2019, n2021, n2025, n2027, n2029, n2031, n2033, n2035, n2037, n2039, n2041, n2043, n1997, n1999, n2003, n2005, n2007, n2009, n2011, n2013;
    wire n2015, n2017, n1983, n1985, n1987, n1989, n1991, n1993, n1995, n2001, n1849, n2096, N869, n1851, n1975, n5816, n1852, n3116, n1853, n1942;
    wire n5849, n2782, n2098, n1935, n2047, n2073, n1969, n2060, n2061, n2069, n2070, n2075, n2076, n2080, n2081, n2044, n2045, n2049, n2050, n2052;
    wire n2053, n2055, n2056, n2083, n2084, n2063, n2064, n2066, n2067, n2089, n2090, n2092, n2093, n5845, n5917, n5782, n2785, n2719, n6064, n6065;
    wire n5996, n5997, n5886, n2591, n2957, n5936, n5789, n1909, n5643, n1910, n5647, n1911, n5649, n1912, n5651, n1913, n5655, n1914, n5657, n1915;
    wire n5665, n1916, n5667, n1917, n5669, n1918, n5671, n1919, n5798, n1920, n5804, n1921, n5866, n1922, n5871, n1923, n5975, n1924, n6012, n1925;
    wire n6032, n1926, n6035, n1927, n6009, n1928, n6081, n1929, n6115, n5780, n6000, n1930, n5844, n5846, n1931, n5890, n5874, n4707, n1932, n6014;
    wire n6061, n4703, n1933, n6039, n5814, n4705, n1934, n5785, n5784, n1937, n5879, n1938, n5946, n1939, n6018, n1940, n6059, n6091, n6090, n1943;
    wire n6107, n1944, n6122, n1945, n5776, n1946, n6019, n1947, n6086, n5763, n1948, n5777, n1949, n6020, n1950, n6044, n1951, n6087, n1952, n6108;
    wire n4663, n1954, n5801, n6067, n1955, n1956, n6071, n5788, n1957, n4692, n1958, n5949, n2892, n1959, n5915, n2953, n1960, n1961, n5865, n5803;
    wire n1962, n5820, n2097, n2115, n1963, n6050, n1964, n1965, n5773, n5783, n1966, n6069, n6021, n1967, n6003, n1968, n5960, n6024, n2714, n1970;
    wire n6080, n6045, n1971, n5799, n2954, n1972, n5756, n2781, n1973, n6073, n6072, n1976, n5812, n5791, n2655, n1977, n5750, n2651, n1978, n5938;
    wire n2715, n2844, n1979, n5830, n2116, n1980, n5847, n1981, n4146, n4145, n4147, n4148, n4173, n4172, n4174, n4175, n4189, n4188, n4190, n4191;
    wire n4205, n4204, n4206, n4207, n4221, n4220, n4222, n4223, n4237, n4236, n4238, n4239, n4253, n4252, n4254, n4255, n4269, n4268, n4270, n4271;
    wire n4285, n4284, n4286, n4287, n4301, n4300, n4302, n4303, n4317, n4316, n4318, n4319, n4333, n4332, n4334, n4335, n4349, n4348, n4350, n4351;
    wire n4365, n4364, n4366, n4367, n4381, n4380, n4382, n4383, n4397, n4396, n4398, n4399, n4413, n4412, n4414, n4415, n4429, n4428, n4430, n4431;
    wire n4447, n4446, n4448, n4449, n4463, n4462, n4464, n4465, n4479, n4478, n4480, n4481, n4495, n4494, n4496, n4497, n4511, n4510, n4512, n4513;
    wire n4527, n4526, n4528, n4529, n4543, n4542, n4544, n4545, n4559, n4558, n4560, n4561, n4575, n4574, n4576, n4577, n4591, n4590, n4592, n4593;
    wire n4607, n4606, n4608, n4609, n4623, n4622, n4624, n4625, n4639, n4638, n4640, n4641, n5744, n5743, n5742, n5759, n5758, n5810, n5809, n5808;
    wire n5825, n5824, n5823, n5835, n5834, n5833, n5851, n5850, n5878, n5877, n5876, n5907, n5906, n5905, n5908, n5909, n5922, n5921, n5920, n5952;
    wire n5951, n5950, n5967, n5966, n5968, n5969, n5978, n5977, n5976, n5995, n5994, n6017, n6016, n6015, n6042, n6041, n6040, n6063, n6062, n6077;
    wire n6076, n6075, n6078, n6079, n6104, n6103, n6102, n6105, n6106, n4655, n4654, n4656, n4657, n5805, n6109, n6083, n6082, n2101, n5781, n5859;
    wire n2102, n4699, n6001, n4711, n2103, n5883, n2104, n6068, n2105, n5904, n2106, n6038, n5885, n2108, n5926, n5779, n5807, n2109, n5755, n2889;
    wire n2110, n5838, n5860, n2111, n5778, n2112, n5914, n5998, n2113, n2114, n5769, n5925, n5889, n2117, n2118, n4154, n2119, n2120, n4152, n2121;
    wire n2122, n4159, n2123, n2124, n4153, n2125, n4718, n3041, n5676, n2126, n3088, n4925, n3087, n2128, n4949, n2129, n5047, n3086, n2130, n5079;
    wire n2131, n5223, n2132, n5427, n2133, n5551, n2134, n2135, n4014, n2136, n3630, n2137, n3246, n4929, n2138, n4951, n2139, n5049, n2140, n5081;
    wire n2141, n5225, n2142, n5429, n3085, n2143, n5555, n2144, n2145, n3886, n2146, n3694, n2147, n3310, n2148, n3628, n2149, n3244, n2150, n4010;
    wire n4939, n2151, n4959, n2152, n5053, n2153, n5083, n2154, n5295, n2155, n5435, n2156, n5557, n2157, n2158, n3822, n2159, n3566, n2160, n3884;
    wire n2161, n3372, n2162, n4008, n2163, n3624, n2164, n3240, n2165, n4070, n2166, n3686, n2167, n3302, n2168, n4911, n2169, n5481, n2170, n5593;
    wire n4953, n2171, n5055, n2172, n5089, n2173, n5297, n2174, n5437, n2175, n5573, n2176, n2177, n3758, n2178, n3374, n2179, n3182, n2180, n3820;
    wire n2181, n3564, n2182, n3308, n2183, n4006, n2184, n3878, n2185, n3622, n2186, n3238, n2187, n4068, n2188, n3684, n2189, n4913, n2190, n4969;
    wire n2191, n5563, n2192, n5603, n4955, n2193, n5095, n2194, n5303, n2195, n5443, n2196, n5577, n2197, n4785, n2198, n2199, n4142, n2200, n3756;
    wire n2201, n3500, n2202, n3180, n2203, n3562, n2204, n3370, n2205, n3816, n2206, n4004, n2207, n3876, n2208, n3620, n2209, n3236, n2210, n4066;
    wire n2211, n3682, n2212, n3298, n2213, n3854, n2214, n3278, n2215, n4933, n2216, n5041, n2217, n5425, n2218, n5567, n2219, n5597, n2220, n5704;
    wire n4961, n2221, n5071, n2222, n5097, n2223, n5325, n2224, n5461, n2225, n5587, n2226, n5710, n2227, n4793, n2228, n2229, n4078, n2230, n3438;
    wire n2231, n4140, n2232, n3692, n2233, n3754, n2234, n3944, n2235, n3496, n2236, n3368, n2237, n3814, n2238, n3300, n2239, n4002, n2240, n3874;
    wire n2241, n3618, n2242, n3234, n2243, n4062, n2244, n3676, n2245, n3548, n2246, n3420, n2247, n3162, n2248, n4114, n2249, n3984, n2250, n3728;
    wire n2251, n3600, n2252, n3790, n2253, n3470, n2254, n3342, n2255, n3214, n2256, n3916, n2257, n4937, n2258, n5197, n2259, n5315, n2260, n5431;
    wire n2261, n5569, n2262, n5702, n2263, n4805, n4715, N646, n2264, n5045, n2265, n5169, n2266, n5327, n2267, n5445, n2268, n5559, n2269, n5718;
    wire n2270, n2271, n3502, n2272, n4076, n2273, n3436, n2274, n4138, n2275, n3178, n2276, n3752, n2277, n3560, n2278, n3942, n2279, n3494, n2280;
    wire n3366, n2281, n3812, n2282, n4000, n2283, n3872, n2284, n3616, n2285, n3232, n2286, n3678, n2287, n3294, n2288, n4060, n2289, n3542, n2290;
    wire n3158, n2291, n4110, n2292, n3918, n2293, n3662, n2294, n3852, n2295, n3724, n2296, n3468, n2297, n3276, n2298, n3338, n2299, n3974, n2300;
    wire n3782, n2301, n3590, n2302, n3398, n2303, n3206, n2304, n4036, n2305, n4915, n2306, n4957, n2307, n5091, n2308, n5199, n2309, n5321, n2310;
    wire n5471, n2311, n5571, n2312, n5599, n2313, n5706, n2314, n4807, n5061, n2315, n5183, n2316, n5329, n2317, n5455, n2318, n5561, n2319, n5692;
    wire n2320, n4823, n2321, n2322, n4012, n2323, n3882, n2324, n3626, n2325, n3498, n2326, n3242, n2327, n4136, n2328, n3750, n2329, n3558, n2330;
    wire n3940, n2331, n3492, n2332, n3364, n2333, n4064, n2334, n3680, n2335, n3296, n2336, n3998, n2337, n3806, n2338, n3614, n2339, n3422, n2340;
    wire n3230, n2341, n3866, n2342, n3160, n2343, n3540, n2344, n4112, n2345, n4046, n2346, n3726, n2347, n3660, n2348, n3340, n2349, n3914, n2350;
    wire n3466, n2351, n3274, n2352, n3972, n2353, n3780, n2354, n3588, n2355, n3396, n2356, n3204, n2357, n3842, n2358, n3136, n2359, n4917, n2360;
    wire n4965, n2361, n5093, n2362, n5211, n2363, n5323, n2364, n5475, n2365, n5575, n2366, n5605, n2367, n5708, n2368, n4809, n5057, n2369, n5185;
    wire n2370, n5305, n2371, n5457, n2372, n5565, n2373, n5698, n2374, n4795, n2375, n4827, n2376, n2377, n4074, n2378, n3818, n2379, n3690, n2380;
    wire n3434, n2381, n3306, n2382, n3176, n2383, n4134, n2384, n3748, n2385, n3938, n2386, n3490, n2387, n3362, n2388, n3870, n2389, n3996, n2390;
    wire n3804, n2391, n3612, n2392, n3228, n2393, n4058, n2394, n3674, n2395, n3546, n2396, n3418, n2397, n3290, n2398, n3156, n2399, n4108, n2400;
    wire n3850, n2401, n3722, n2402, n3912, n2403, n3464, n2404, n3336, n2405, n3970, n2406, n3778, n2407, n3650, n2408, n3522, n2409, n3394, n2410;
    wire n3202, n2411, n4032, n2412, n3584, n2413, n3264, n2414, n3134, n2415, n4919, n2416, n5043, n2417, n5167, n2418, n5213, n2419, n5335, n2420;
    wire n5479, n2421, n5581, n2422, n5712, n2423, n4811, n2424, n5827, n4963, n2425, n5067, n2426, n5191, n2427, n5307, n2428, n5463, n2429, n5589;
    wire n2430, n5724, n2431, n4831, n2432, n2433, n4072, n2434, n3880, n2435, n3688, n2436, n3432, n2437, n3304, n2438, n3174, n2439, n4132, n2440;
    wire n3746, n2441, n3936, n2442, n3488, n2443, n3360, n2444, n3994, n2445, n3802, n2446, n3610, n2447, n3226, n2448, n3864, n2449, n3672, n2450;
    wire n3544, n2451, n3416, n2452, n3288, n2453, n4054, n2454, n3154, n2455, n4106, n2456, n3720, n2457, n3910, n2458, n3462, n2459, n3334, n2460;
    wire n4034, n2461, n3586, n2462, n3266, n2463, n3968, n2464, n3776, n2465, n3648, n2466, n3520, n2467, n3392, n2468, n3200, n2469, n3838, n2470;
    wire n3132, n2471, n5069, n2472, n5171, n2473, n5215, n2474, n5337, n2475, n5433, n2476, n5680, n2477, n5732, n2478, n4813, n2479, n5963, n2481;
    wire n5928, n5930, n5931, n5932, n4967, n2482, n5201, n2483, n5311, n2484, n5465, n2485, n5595, n2486, n5700, n2487, n4835, n2488, n2489, n3430;
    wire n2490, n3556, n2491, n3172, n2492, n4130, n2493, n3744, n2494, n3934, n2495, n3486, n2496, n3358, n2497, n4056, n2498, n3800, n2499, n3608;
    wire n2500, n3224, n2501, n3990, n2502, n3862, n2503, n3670, n2504, n3414, n2505, n3286, n2506, n3538, n2507, n3152, n2508, n3460, n2509, n3840;
    wire n2510, n4094, n2511, n3966, n2512, n3774, n2513, n3646, n2514, n3518, n2515, n3326, n2516, n3198, n2517, n4028, n2518, n3900, n2519, n3708;
    wire n2520, n3580, n2521, n3388, n2522, n3260, n2523, n3130, n2524, n4921, n2525, n5051, n2526, n5175, n2527, n5217, n2528, n5339, n2529, n5447;
    wire n2530, n5553, n2531, n5714, n2532, n4787, n2533, n4815, n2534, n5990, n5852, n5855, n5856, n2535, n2536, n2538, n5940, n5942, n5943, n5944;
    wire n5037, N710, n2539, n5075, n2540, n5203, n2541, n5317, n2542, n5467, n2543, n5684, n2544, n5726, n2545, n4841, n2546, n2547, n3428, n2548;
    wire n3810, n2549, n3554, n2550, n3170, n2551, n3484, n2552, n3992, n2553, n3926, n2554, n3734, n2555, n3606, n2556, n3350, n2557, n3222, n2558;
    wire n4116, n2559, n3860, n2560, n3668, n2561, n3412, n2562, n3284, n2563, n4050, n2564, n3536, n2565, n3150, n2566, n3788, n2567, n3458, n2568;
    wire n4030, n2569, n3902, n2570, n3710, n2571, n3582, n2572, n3390, n2573, n3262, n2574, n4092, n2575, n3964, n2576, n3836, n2577, n3644, n2578;
    wire n3516, n2579, n3324, n2580, n3196, n2581, n3768, n2582, n4927, n2583, n5059, n2584, n5179, n2585, n5219, n2586, n5341, n2587, n5449, n2588;
    wire n5607, n2589, n5734, n2590, n4817, n6074, n5899, n2592, n2593, n2594, n5039, n2596, n5173, n2597, n5331, n2598, n5469, n2599, n5601, n2600;
    wire n4837, n2601, n2602, n3950, n2603, n3426, n2604, n3552, n2605, n3168, n2606, n3482, n2607, n4118, n2608, n3798, n2609, n4052, n2610, n3924;
    wire n2611, n3732, n2612, n3604, n2613, n3348, n2614, n3220, n2615, n3986, n2616, n3858, n2617, n3666, n2618, n3410, n2619, n3282, n2620, n3534;
    wire n2621, n3148, n2622, n3456, n2623, n3772, n2624, n4090, n2625, n3962, n2626, n3834, n2627, n3642, n2628, n3514, n2629, n3322, n2630, n3194;
    wire n2631, n4024, n2632, n3896, n2633, n3704, n2634, n3576, n2635, n3384, n2636, n3256, n2637, n3128, n3112, n3094, n2638, n2639, n4943, n2640;
    wire n5063, n2641, n5181, n2642, n5221, n2643, n5349, n2644, n5451, n2645, n5686, n2646, n5716, n2647, n4782, n2648, n4819, n2650, n5985, n5987;
    wire n5988, n5989, n5822, n5792, n2652, n5819, n2784, n2653, n2654, n5875, n5754, n2656, n5077, n2658, n5205, n2659, n5319, n2660, n5473, n2661;
    wire n5609, n2662, n4799, n2663, n2664, n3948, n2665, n4128, n2666, n3808, n2667, n3424, n2668, n3550, n2669, n3166, n2670, n3480, n2671, n3988;
    wire n2672, n3922, n2673, n3730, n2674, n3602, n2675, n3346, n2676, n3218, n2677, n4048, n2678, n3856, n2679, n3664, n2680, n3408, n2681, n3280;
    wire n2682, n3532, n2683, n3786, n2684, n3146, n2685, n4104, n2686, n3454, n2687, n4026, n2688, n3898, n2689, n3706, n2690, n3578, n2691, n3386;
    wire n2692, n3258, n2693, n4088, n2694, n3960, n2695, n3832, n2696, n3640, n2697, n3512, n2698, n3320, n2699, n3192, n2700, n3766, n3110, n2701;
    wire n2702, n5065, n2703, n5187, n2704, n5299, n2705, n5343, n2706, n5439, n2707, n5579, n2708, n5688, n2709, n5722, n2710, n4789, n2711, n4825;
    wire n5840, n6002, n5903, n2713, n5972, n5934, n2716, n5757, n6117, n5916, n4701, n4931, n2721, n5207, n2722, n5333, n2723, n5477, n2724, n5678;
    wire N614, n2725, n4803, n2726, n2727, n3946, n2728, n4126, n2729, n3742, n2730, n3868, n2731, n3356, n2732, n3478, n2733, n3796, n2734, n3920;
    wire n2735, n3982, n2736, n3598, n2737, n3406, n2738, n4044, n2739, n3212, n2740, n3658, n2741, n3530, n2742, n3272, n2743, n3144, n2744, n4102;
    wire n2745, n3718, n2746, n3332, n2747, n3452, n2748, n3770, n2749, n4022, n2750, n3894, n2751, n3638, n2752, n3510, n2753, n3382, n2754, n3254;
    wire n2755, n3126, n2756, n4084, n2757, n3956, n2758, n3828, n2759, n3700, n2760, n3572, n2761, n3444, n2762, n3316, n2763, n3188, n3108, n2764;
    wire n2765, n4945, n2766, n5073, n2767, n5189, n2768, n5301, n2769, n5353, n2770, n5453, n2771, n5583, n2772, n5694, n2773, n5720, n2774, n4791;
    wire n2775, n4829, n2776, n3104, n6089, n2778, n6094, n6095, n6096, n2780, n5772, n5209, n2786, n5345, n2787, n5682, n2788, n5739, n2789, n4821;
    wire n2790, n2791, n4124, n2792, n3932, n2793, n3740, n2794, n3292, n2795, n3164, n2796, n3476, n2797, n3794, n2798, n3344, n2799, n3216, n2800;
    wire n3980, n2801, n3596, n2802, n3404, n2803, n4042, n2804, n3848, n2805, n3656, n2806, n3528, n2807, n3142, n2808, n4100, n2809, n3908, n2810;
    wire n3716, n2811, n3450, n2812, n4086, n2813, n3958, n2814, n3830, n2815, n3702, n2816, n3574, n2817, n3446, n2818, n3318, n2819, n3190, n2820;
    wire n4020, n2821, n3892, n2822, n3764, n2823, n3636, n2824, n3508, n2825, n3380, n2826, n3252, n2827, n3124, n2828, n4947, n2829, n5085, n2830;
    wire n5193, n2831, n5309, n2832, n5423, n2833, n5459, n2834, n5585, n2835, n5690, n2836, n5730, n2837, n4797, n2838, n4833, n4971, n2839, n3096;
    wire n3099, n2840, n3097, n2841, n5831, n2842, n5918, n2843, n2846, n6118, n2848, n4700, n2850, n4122, n2851, n3930, n2852, n3738, n2853, n3354;
    wire n2854, n3474, n2855, n3978, n2856, n3594, n2857, n3402, n2858, n3210, n2859, n4040, n2860, n3784, n2861, n3846, n2862, n3654, n2863, n3526;
    wire n2864, n3270, n2865, n3140, n2866, n4098, n2867, n3906, n2868, n3714, n2869, n3330, n2870, n4018, n2871, n3890, n2872, n3762, n2873, n3634;
    wire n2874, n3506, n2875, n3378, n2876, n3250, n2877, n3122, n2878, n4080, n2879, n3952, n2880, n3824, n2881, n3696, n2882, n3568, n2883, n3440;
    wire n2884, n3312, n2885, n3184, n3114, n2886, n2887, n4696, n2888, n4445, n4144, n2895, n4941, n2896, n5177, n2897, n5728, n2898, n2899, n4120;
    wire n2900, n3928, n2901, n3736, n2902, n3352, n2903, n3792, n2904, n3472, n2905, n3976, n2906, n3592, n2907, n3400, n2908, n3208, n2909, n4038;
    wire n2910, n3844, n2911, n3652, n2912, n3524, n2913, n3268, n2914, n3138, n2915, n4096, n2916, n3904, n2917, n3712, n2918, n3328, n2919, n3448;
    wire n2920, n4082, n2921, n3954, n2922, n3826, n2923, n3698, n2924, n3570, n2925, n3442, n2926, n3314, n2927, n3186, n2928, n4016, n2929, n3888;
    wire n2930, n3760, n2931, n3632, n2932, n3504, n2933, n3376, n2934, n3248, n2935, n3119, n2936, n5087, n2937, n5195, n2938, n5313, n2939, n5347;
    wire n2940, n5441, n2941, n5591, n2942, n5696, n2943, n5736, n2944, n4801, n2945, n4839, n5227, n2946, n5355, n2947, n5483, n2948, n5741, n2949;
    wire n2980, n2950, n5737, n2952, n2956, n3098, n3113, n4168, n3089, n3062, n3081, n3055, n3059, n3053, n3061, n3054, n3058, n3063, n3060, n3057;
    wire n3056, n3052, n3051, n3078, n3070, n3075, n3067, n3080, n3072, n3064, n3077, n3069, n3074, n3066, n3079, n3076, n3073, n3071, n3068, n3065;
    wire n3009, n3012, n3001, n2993, n3006, n2998, n2990, n3011, n3003, n2995, n2987, n3008, n3000, n2992, n3005, n2997, n2989, n3010, n3007, n3004;
    wire n3002, n2999, n2996, n2994, n2991, n2988, n2986, n2985, n2982, n2984, n2981, n2983, n2977, n2979, n2978, n3016, n3049, n3015, n3027, n3032;
    wire n3039, n3017, n3022, n3038, n3025, n3030, n3042, n3035, n3020, n3028, n3033, n3018, n3040, n3023, n3037, n3026, n3029, n3031, n3034, n3019;
    wire n3021, n3024, n3036, n3045, n3043, n3044, n3046, n3047, n3048, n3093, n3092, n3120, n3083, n3084, n3082, n3013, n3014, n3050, N902, N934;
    wire n3091, n2976, n3090, N1029, N870, w_mem_inst_N640, w_mem_inst_N672, n3117, N997, w_mem_inst_N639, w_mem_inst_N607, N837, N1579, N1547, N774, N742, N678, N582, N550, n3095;
    wire n3101, n3102, n3105, n3106, n3107, n3109, n3111, n3118, n3121, n3123, n3125, n3127, n3129, n3131, n3133, n3135, n3137, n3139, n3141, n3143;
    wire n3145, n3147, n3149, n3151, n3153, n3155, n3157, n3159, n3161, n3163, n3165, n3167, n3169, n3171, n3173, n3175, n3177, n3179, n3181, n3183;
    wire n3185, n3187, n3189, n3191, n3193, n3195, n3197, n3199, n3201, n3203, n3205, n3207, n3209, n3211, n3213, n3215, n3217, n3219, n3221, n3223;
    wire n3225, n3227, n3229, n3231, n3233, n3235, n3237, n3239, n3241, n3243, n3245, n3247, n3249, n3251, n3253, n3255, n3257, n3259, n3261, n3263;
    wire n3265, n3267, n3269, n3271, n3273, n3275, n3277, n3279, n3281, n3283, n3285, n3287, n3289, n3291, n3293, n3295, n3297, n3299, n3301, n3303;
    wire n3305, n3307, n3309, n3311, n3313, n3315, n3317, n3319, n3321, n3323, n3325, n3327, n3329, n3331, n3333, n3335, n3337, n3339, n3341, n3343;
    wire n3345, n3347, n3349, n3351, n3353, n3355, n3357, n3359, n3361, n3363, n3365, n3367, n3369, n3371, n3373, n3375, n3377, n3379, n3381, n3383;
    wire n3385, n3387, n3389, n3391, n3393, n3395, n3397, n3399, n3401, n3403, n3405, n3407, n3409, n3411, n3413, n3415, n3417, n3419, n3421, n3423;
    wire n3425, n3427, n3429, n3431, n3433, n3435, n3437, n3439, n3441, n3443, n3445, n3447, n3449, n3451, n3453, n3455, n3457, n3459, n3461, n3463;
    wire n3465, n3467, n3469, n3471, n3473, n3475, n3477, n3479, n3481, n3483, n3485, n3487, n3489, n3491, n3493, n3495, n3497, n3499, n3501, n3503;
    wire n3505, n3507, n3509, n3511, n3513, n3515, n3517, n3519, n3521, n3523, n3525, n3527, n3529, n3531, n3533, n3535, n3537, n3539, n3541, n3543;
    wire n3545, n3547, n3549, n3551, n3553, n3555, n3557, n3559, n3561, n3563, n3565, n3567, n3569, n3571, n3573, n3575, n3577, n3579, n3581, n3583;
    wire n3585, n3587, n3589, n3591, n3593, n3595, n3597, n3599, n3601, n3603, n3605, n3607, n3609, n3611, n3613, n3615, n3617, n3619, n3621, n3623;
    wire n3625, n3627, n3629, n3631, n3633, n3635, n3637, n3639, n3641, n3643, n3645, n3647, n3649, n3651, n3653, n3655, n3657, n3659, n3661, n3663;
    wire n3665, n3667, n3669, n3671, n3673, n3675, n3677, n3679, n3681, n3683, n3685, n3687, n3689, n3691, n3693, n3695, n3697, n3699, n3701, n3703;
    wire n3705, n3707, n3709, n3711, n3713, n3715, n3717, n3719, n3721, n3723, n3725, n3727, n3729, n3731, n3733, n3735, n3737, n3739, n3741, n3743;
    wire n3745, n3747, n3749, n3751, n3753, n3755, n3757, n3759, n3761, n3763, n3765, n3767, n3769, n3771, n3773, n3775, n3777, n3779, n3781, n3783;
    wire n3785, n3787, n3789, n3791, n3793, n3795, n3797, n3799, n3801, n3803, n3805, n3807, n3809, n3811, n3813, n3815, n3817, n3819, n3821, n3823;
    wire n3825, n3827, n3829, n3831, n3833, n3835, n3837, n3839, n3841, n3843, n3845, n3847, n3849, n3851, n3853, n3855, n3857, n3859, n3861, n3863;
    wire n3865, n3867, n3869, n3871, n3873, n3875, n3877, n3879, n3881, n3883, n3885, n3887, n3889, n3891, n3893, n3895, n3897, n3899, n3901, n3903;
    wire n3905, n3907, n3909, n3911, n3913, n3915, n3917, n3919, n3921, n3923, n3925, n3927, n3929, n3931, n3933, n3935, n3937, n3939, n3941, n3943;
    wire n3945, n3947, n3949, n3951, n3953, n3955, n3957, n3959, n3961, n3963, n3965, n3967, n3969, n3971, n3973, n3975, n3977, n3979, n3981, n3983;
    wire n3985, n3987, n3989, n3991, n3993, n3995, n3997, n3999, n4001, n4003, n4005, n4007, n4009, n4011, n4013, n4015, n4017, n4019, n4021, n4023;
    wire n4025, n4027, n4029, n4031, n4033, n4035, n4037, n4039, n4041, n4043, n4045, n4047, n4049, n4051, n4053, n4055, n4057, n4059, n4061, n4063;
    wire n4065, n4067, n4069, n4071, n4073, n4075, n4077, n4079, n4081, n4083, n4085, n4087, n4089, n4091, n4093, n4095, n4097, n4099, n4101, n4103;
    wire n4105, n4107, n4109, n4111, n4113, n4115, n4117, n4119, n4121, n4123, n4125, n4127, n4129, n4131, n4133, n4135, n4137, n4139, n4141, n4143;
    wire n4149, n4150, n4151, n4155, n4156, n4157, n4158, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4171, n4176, n4177, n4178, n4179;
    wire n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203;
    wire n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231;
    wire n4232, n4233, n4234, n4235, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4256, n4257, n4258, n4259;
    wire n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283;
    wire n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311;
    wire n4312, n4313, n4314, n4315, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4336, n4337, n4338, n4339;
    wire n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363;
    wire n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391;
    wire n4392, n4393, n4394, n4395, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4416, n4417, n4418, n4419;
    wire n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4443, n4444;
    wire n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473;
    wire n4474, n4475, n4476, n4477, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4498, n4499, n4500, n4501;
    wire n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525;
    wire n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553;
    wire n4554, n4555, n4556, n4557, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4578, n4579, n4580, n4581;
    wire n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605;
    wire n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633;
    wire n4634, n4635, n4636, n4637, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4658, n4659, n4660, n4661;
    wire n4662, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682;
    wire n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4693, n4694, n4695, n4697, n4698, n4702, n4704, n4706, n4708, n4709, n4710;
    wire n4712, n4714, n4716, n4717, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734;
    wire n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754;
    wire n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774;
    wire n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4784, n4786, n4788, n4790, n4792, n4794, n4796, n4798, n4800, n4802, n4804, n4806, n4808;
    wire n4810, n4812, n4814, n4816, n4818, n4820, n4822, n4824, n4826, n4828, n4830, n4832, n4834, n4836, n4838, n4840, n4842, n4843, n4844, n4845;
    wire n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865;
    wire n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885;
    wire n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905;
    wire n4906, n4907, n4908, n4909, n4910, n4912, n4914, n4916, n4918, n4920, n4922, n4923, n4924, n4926, n4928, n4930, n4932, n4934, n4935, n4936;
    wire n4938, n4940, n4942, n4944, n4946, n4948, n4950, n4952, n4954, n4956, n4958, n4960, n4962, n4964, n4966, n4968, n4970, n4972, n4973, n4974;
    wire n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994;
    wire n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014;
    wire n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034;
    wire n5035, n5036, n5038, n5040, n5042, n5044, n5046, n5048, n5050, n5052, n5054, n5056, n5058, n5060, n5062, n5064, n5066, n5068, n5070, n5072;
    wire n5074, n5076, n5078, n5080, n5082, n5084, n5086, n5088, n5090, n5092, n5094, n5096, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105;
    wire n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125;
    wire n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145;
    wire n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165;
    wire n5166, n5168, n5170, n5172, n5174, n5176, n5178, n5180, n5182, n5184, n5186, n5188, n5190, n5192, n5194, n5196, n5198, n5200, n5202, n5204;
    wire n5206, n5208, n5210, n5212, n5214, n5216, n5218, n5220, n5222, n5224, n5226, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236;
    wire n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256;
    wire n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276;
    wire n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5296, n5298;
    wire n5300, n5302, n5304, n5306, n5308, n5310, n5312, n5314, n5316, n5318, n5320, n5322, n5324, n5326, n5328, n5330, n5332, n5334, n5336, n5338;
    wire n5340, n5342, n5344, n5346, n5348, n5350, n5351, n5352, n5354, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366;
    wire n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386;
    wire n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406;
    wire n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5424, n5426, n5428, n5430;
    wire n5432, n5434, n5436, n5438, n5440, n5442, n5444, n5446, n5448, n5450, n5452, n5454, n5456, n5458, n5460, n5462, n5464, n5466, n5468, n5470;
    wire n5472, n5474, n5476, n5478, n5480, n5482, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497;
    wire n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517;
    wire n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537;
    wire n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5552, n5554, n5556, n5558, n5560, n5562, n5564;
    wire n5566, n5568, n5570, n5572, n5574, n5576, n5578, n5580, n5582, n5584, n5586, n5588, n5590, n5592, n5594, n5596, n5598, n5600, n5602, n5604;
    wire n5606, n5608, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627;
    wire n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5644, n5645, n5646, n5648, n5650;
    wire n5652, n5653, n5654, n5656, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5666, n5668, n5670, n5672, n5673, n5674, n5675, n5677, n5679;
    wire n5681, n5683, n5685, n5687, n5689, n5691, n5693, n5695, n5697, n5699, n5701, n5703, n5705, n5707, n5709, n5711, n5713, n5715, n5717, n5719;
    wire n5721, n5723, n5725, n5727, n5729, n5731, n5733, n5735, n5738, n5740, n5745, n5746, n5747, n5748, n5753, n5760, n5761, n5762, n5764, n5765;
    wire n5766, n5767, n5768, n5774, n5775, n5787, n5790, n5794, n5795, n5796, n5797, n5800, n5802, n5806, n5811, n5813, n5815, n5817, n5818, n5826;
    wire n5828, n5829, n5832, n5836, n5841, n5842, n5854, n5857, n5858, n5862, n5863, n5864, n5868, n5869, n5870, n5872, n5873, n5880, n5881, n5882;
    wire n5884, n5887, n5888, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5900, n5901, n5902, n5910, n5911, n5913, n5919, n5923, n5924;
    wire n5927, n5929, n5933, n5935, n5937, n5939, n5941, n5945, n5947, n5948, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5961, n5962, n5964;
    wire n5965, n5970, n5973, n5974, n5979, n5980, n5982, n5983, n5984, n5986, n5992, n5993, n5999, n6004, n6005, n6006, n6007, n6008, n6010, n6011;
    wire n6013, n6022, n6023, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6034, n6036, n6037, n6043, n6046, n6047, n6048, n6049, n6051, n6052;
    wire n6053, n6054, n6055, n6056, n6057, n6058, n6060, n6066, n6070, n6084, n6085, n6088, n6092, n6093, n6097, n6098, n6099, n6100, n6101, n6110;
    wire n6111, n6112, n6113, n6114, n6116, n6119, n6120, n6121, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134;
    wire n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154;
    wire n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174;
    wire n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, puf_0_wire_0;
    wire puf_0_wire_1, puf_0_wire_2, puf_0_wire_3, puf_1_wire_0, puf_1_wire_1, puf_1_wire_2, puf_1_wire_3, puf_2_wire_0, puf_2_wire_1, puf_2_wire_2, puf_2_wire_3, puf_3_wire_0, puf_3_wire_1, puf_3_wire_2, puf_3_wire_3, puf_4_wire_0, puf_4_wire_1, puf_4_wire_2, puf_4_wire_3, puf_5_wire_0;
    wire puf_5_wire_1, puf_5_wire_2, puf_5_wire_3, puf_6_wire_0, puf_6_wire_1, puf_6_wire_2, puf_6_wire_3, puf_7_wire_0, puf_7_wire_1, puf_7_wire_2, puf_7_wire_3, puf_8_wire_0, puf_8_wire_1, puf_8_wire_2, puf_8_wire_3, puf_9_wire_0, puf_9_wire_1, puf_9_wire_2, puf_9_wire_3, puf_10_wire_0;
    wire puf_10_wire_1, puf_10_wire_2, puf_10_wire_3, puf_11_wire_0, puf_11_wire_1, puf_11_wire_2, puf_11_wire_3, puf_12_wire_0, puf_12_wire_1, puf_12_wire_2, puf_12_wire_3, puf_13_wire_0, puf_13_wire_1, puf_13_wire_2, puf_13_wire_3, puf_14_wire_0, puf_14_wire_1, puf_14_wire_2, puf_14_wire_3, puf_15_wire_0;
    wire puf_15_wire_1, puf_15_wire_2, puf_15_wire_3;
    wire [1:0] sha256_ctrl_reg;
    wire [5:0] t_ctr_reg;
    wire [31:0] d_reg;
    wire [31:0] e_reg;
    wire [31:0] f_reg;
    wire [31:0] g_reg;
    wire [31:0] h_reg;
    wire [31:0] a_reg;
    wire [31:0] b_reg;
    wire [31:0] c_reg;
    wire [511:0] w_mem_inst_w_mem;
    wire [5:0] w_mem_inst_w_ctr_reg;
    wire [31:2] w_mem_inst_add_2_root_add_945_3_carry;
    wire [31:2] w_mem_inst_add_1_root_add_945_3_carry;
    wire [31:2] w_mem_inst_add_0_root_add_945_3_carry;
    wire [31:0] w_mem_inst_w_new;
    wire [5:2] w_mem_inst_add_1008_carry;
    wire [5:2] add_420_carry;
    wire [31:2] add_392_carry;
    wire [31:0] t1;
    wire [31:2] add_0_root_add_388_carry;
    wire [31:0] t2;
    wire [31:2] add_1_root_add_388_carry;
    wire [31:2] add_0_root_add_317_4_carry;
    wire [31:2] add_1_root_add_317_4_carry;
    wire [30:0] k_data;
    wire [31:2] add_2_root_add_317_4_carry;
    wire [31:2] add_3_root_add_317_4_carry;
    wire [31:2] add_295_carry;
    wire [31:2] add_294_carry;
    wire [31:2] add_293_carry;
    wire [31:2] add_292_carry;
    wire [31:2] add_291_carry;
    wire [31:2] add_290_carry;
    wire [31:2] add_289_carry;
    wire [31:2] add_288_carry;


   DFFPOSX1 sha256_ctrl_reg_reg_0_ ( .CLK(clk),  .D(n1755), .Q(sha256_ctrl_reg[0]));
   DFFPOSX1 t_ctr_reg_reg_5_ ( .CLK(clk),  .D(n1747), .Q(t_ctr_reg[5]));
   DFFPOSX1 sha256_ctrl_reg_reg_1_ ( .CLK(clk),  .D(n1754), .Q(sha256_ctrl_reg[1]));
   DFFPOSX1 t_ctr_reg_reg_0_ ( .CLK(clk),  .D(n1752), .Q(t_ctr_reg[0]));
   DFFPOSX1 t_ctr_reg_reg_1_ ( .CLK(clk),  .D(n1751), .Q(t_ctr_reg[1]));
   DFFPOSX1 t_ctr_reg_reg_2_ ( .CLK(clk),  .D(n1750), .Q(t_ctr_reg[2]));
   DFFPOSX1 t_ctr_reg_reg_3_ ( .CLK(clk),  .D(n1749), .Q(t_ctr_reg[3]));
   DFFPOSX1 t_ctr_reg_reg_4_ ( .CLK(clk),  .D(n1748), .Q(t_ctr_reg[4]));
   DFFPOSX1 digest_valid_reg_reg ( .CLK(clk),  .D(n1753), .Q(digest_valid));
   DFFPOSX1 H3_reg_reg_0_ ( .CLK(clk),  .D(n1746), .Q(digest[128]));
   DFFPOSX1 d_reg_reg_0_ ( .CLK(clk),  .D(n1745), .Q(d_reg[0]));
   DFFPOSX1 e_reg_reg_31_ ( .CLK(clk),  .D(n1651), .Q(e_reg[31]));
   DFFPOSX1 H4_reg_reg_0_ ( .CLK(clk),  .D(n1650), .Q(digest[96]));
   DFFPOSX1 e_reg_reg_0_ ( .CLK(clk),  .D(n1682), .Q(e_reg[0]));
   DFFPOSX1 H4_reg_reg_1_ ( .CLK(clk),  .D(n1649), .Q(digest[97]));
   DFFPOSX1 e_reg_reg_1_ ( .CLK(clk),  .D(n1681), .Q(e_reg[1]));
   DFFPOSX1 H4_reg_reg_2_ ( .CLK(clk),  .D(n1648), .Q(digest[98]));
   DFFPOSX1 e_reg_reg_2_ ( .CLK(clk),  .D(n1680), .Q(e_reg[2]));
   DFFPOSX1 H4_reg_reg_3_ ( .CLK(clk),  .D(n1647), .Q(digest[99]));
   DFFPOSX1 e_reg_reg_3_ ( .CLK(clk),  .D(n1679), .Q(e_reg[3]));
   DFFPOSX1 H4_reg_reg_4_ ( .CLK(clk),  .D(n1646), .Q(digest[100]));
   DFFPOSX1 e_reg_reg_4_ ( .CLK(clk),  .D(n1678), .Q(e_reg[4]));
   DFFPOSX1 H4_reg_reg_5_ ( .CLK(clk),  .D(n1645), .Q(digest[101]));
   DFFPOSX1 e_reg_reg_5_ ( .CLK(clk),  .D(n1677), .Q(e_reg[5]));
   DFFPOSX1 H4_reg_reg_6_ ( .CLK(clk),  .D(n1644), .Q(digest[102]));
   DFFPOSX1 e_reg_reg_6_ ( .CLK(clk),  .D(n1676), .Q(e_reg[6]));
   DFFPOSX1 H4_reg_reg_7_ ( .CLK(clk),  .D(n1643), .Q(digest[103]));
   DFFPOSX1 e_reg_reg_7_ ( .CLK(clk),  .D(n1675), .Q(e_reg[7]));
   DFFPOSX1 H4_reg_reg_8_ ( .CLK(clk),  .D(n1642), .Q(digest[104]));
   DFFPOSX1 e_reg_reg_8_ ( .CLK(clk),  .D(n1674), .Q(e_reg[8]));
   DFFPOSX1 H4_reg_reg_9_ ( .CLK(clk),  .D(n1641), .Q(digest[105]));
   DFFPOSX1 e_reg_reg_9_ ( .CLK(clk),  .D(n1673), .Q(e_reg[9]));
   DFFPOSX1 H4_reg_reg_10_ ( .CLK(clk),  .D(n1640), .Q(digest[106]));
   DFFPOSX1 e_reg_reg_10_ ( .CLK(clk),  .D(n1672), .Q(e_reg[10]));
   DFFPOSX1 H4_reg_reg_11_ ( .CLK(clk),  .D(n1639), .Q(digest[107]));
   DFFPOSX1 e_reg_reg_11_ ( .CLK(clk),  .D(n1671), .Q(e_reg[11]));
   DFFPOSX1 H4_reg_reg_12_ ( .CLK(clk),  .D(n1638), .Q(digest[108]));
   DFFPOSX1 e_reg_reg_12_ ( .CLK(clk),  .D(n1670), .Q(e_reg[12]));
   DFFPOSX1 H4_reg_reg_13_ ( .CLK(clk),  .D(n1637), .Q(digest[109]));
   DFFPOSX1 e_reg_reg_13_ ( .CLK(clk),  .D(n1669), .Q(e_reg[13]));
   DFFPOSX1 H4_reg_reg_14_ ( .CLK(clk),  .D(n1636), .Q(digest[110]));
   DFFPOSX1 e_reg_reg_14_ ( .CLK(clk),  .D(n1668), .Q(e_reg[14]));
   DFFPOSX1 H4_reg_reg_15_ ( .CLK(clk),  .D(n1635), .Q(digest[111]));
   DFFPOSX1 e_reg_reg_15_ ( .CLK(clk),  .D(n1667), .Q(e_reg[15]));
   DFFPOSX1 H4_reg_reg_16_ ( .CLK(clk),  .D(n1634), .Q(puf_0_wire_3));
   DFFPOSX1 e_reg_reg_16_ ( .CLK(clk),  .D(n1666), .Q(e_reg[16]));
   DFFPOSX1 H4_reg_reg_17_ ( .CLK(clk),  .D(n1633), .Q(digest[113]));
   DFFPOSX1 e_reg_reg_17_ ( .CLK(clk),  .D(n1665), .Q(e_reg[17]));
   DFFPOSX1 H4_reg_reg_18_ ( .CLK(clk),  .D(n1632), .Q(digest[114]));
   DFFPOSX1 e_reg_reg_18_ ( .CLK(clk),  .D(n1664), .Q(e_reg[18]));
   DFFPOSX1 H4_reg_reg_19_ ( .CLK(clk),  .D(n1631), .Q(digest[115]));
   DFFPOSX1 e_reg_reg_19_ ( .CLK(clk),  .D(n1663), .Q(e_reg[19]));
   DFFPOSX1 H4_reg_reg_20_ ( .CLK(clk),  .D(n1630), .Q(digest[116]));
   DFFPOSX1 e_reg_reg_20_ ( .CLK(clk),  .D(n1662), .Q(e_reg[20]));
   DFFPOSX1 H4_reg_reg_21_ ( .CLK(clk),  .D(n1629), .Q(digest[117]));
   DFFPOSX1 e_reg_reg_21_ ( .CLK(clk),  .D(n1661), .Q(e_reg[21]));
   DFFPOSX1 H4_reg_reg_22_ ( .CLK(clk),  .D(n1628), .Q(digest[118]));
   DFFPOSX1 e_reg_reg_22_ ( .CLK(clk),  .D(n1660), .Q(e_reg[22]));
   DFFPOSX1 H4_reg_reg_23_ ( .CLK(clk),  .D(n1627), .Q(digest[119]));
   DFFPOSX1 e_reg_reg_23_ ( .CLK(clk),  .D(n1659), .Q(e_reg[23]));
   DFFPOSX1 H4_reg_reg_24_ ( .CLK(clk),  .D(n1626), .Q(digest[120]));
   DFFPOSX1 e_reg_reg_24_ ( .CLK(clk),  .D(n1658), .Q(e_reg[24]));
   DFFPOSX1 H4_reg_reg_25_ ( .CLK(clk),  .D(n1625), .Q(digest[121]));
   DFFPOSX1 e_reg_reg_25_ ( .CLK(clk),  .D(n1657), .Q(e_reg[25]));
   DFFPOSX1 H4_reg_reg_26_ ( .CLK(clk),  .D(n1624), .Q(digest[122]));
   DFFPOSX1 e_reg_reg_26_ ( .CLK(clk),  .D(n1656), .Q(e_reg[26]));
   DFFPOSX1 H4_reg_reg_27_ ( .CLK(clk),  .D(n1623), .Q(digest[123]));
   DFFPOSX1 e_reg_reg_27_ ( .CLK(clk),  .D(n1655), .Q(e_reg[27]));
   DFFPOSX1 H4_reg_reg_28_ ( .CLK(clk),  .D(n1622), .Q(digest[124]));
   DFFPOSX1 e_reg_reg_28_ ( .CLK(clk),  .D(n1654), .Q(e_reg[28]));
   DFFPOSX1 H4_reg_reg_29_ ( .CLK(clk),  .D(n1621), .Q(digest[125]));
   DFFPOSX1 e_reg_reg_29_ ( .CLK(clk),  .D(n1653), .Q(e_reg[29]));
   DFFPOSX1 H4_reg_reg_30_ ( .CLK(clk),  .D(n1620), .Q(digest[126]));
   DFFPOSX1 e_reg_reg_30_ ( .CLK(clk),  .D(n1652), .Q(e_reg[30]));
   DFFPOSX1 H4_reg_reg_31_ ( .CLK(clk),  .D(n1619), .Q(digest[127]));
   DFFPOSX1 f_reg_reg_31_ ( .CLK(clk),  .D(n1587), .Q(f_reg[31]));
   DFFPOSX1 H5_reg_reg_0_ ( .CLK(clk),  .D(n1586), .Q(digest[64]));
   DFFPOSX1 f_reg_reg_0_ ( .CLK(clk),  .D(n1618), .Q(f_reg[0]));
   DFFPOSX1 H5_reg_reg_1_ ( .CLK(clk),  .D(n1585), .Q(digest[65]));
   DFFPOSX1 f_reg_reg_1_ ( .CLK(clk),  .D(n1617), .Q(f_reg[1]));
   DFFPOSX1 H5_reg_reg_2_ ( .CLK(clk),  .D(n1584), .Q(digest[66]));
   DFFPOSX1 f_reg_reg_2_ ( .CLK(clk),  .D(n1616), .Q(f_reg[2]));
   DFFPOSX1 H5_reg_reg_3_ ( .CLK(clk),  .D(n1583), .Q(digest[67]));
   DFFPOSX1 f_reg_reg_3_ ( .CLK(clk),  .D(n1615), .Q(f_reg[3]));
   DFFPOSX1 H5_reg_reg_4_ ( .CLK(clk),  .D(n1582), .Q(digest[68]));
   DFFPOSX1 f_reg_reg_4_ ( .CLK(clk),  .D(n1614), .Q(f_reg[4]));
   DFFPOSX1 H5_reg_reg_5_ ( .CLK(clk),  .D(n1581), .Q(digest[69]));
   DFFPOSX1 f_reg_reg_5_ ( .CLK(clk),  .D(n1613), .Q(f_reg[5]));
   DFFPOSX1 H5_reg_reg_6_ ( .CLK(clk),  .D(n1580), .Q(digest[70]));
   DFFPOSX1 f_reg_reg_6_ ( .CLK(clk),  .D(n1612), .Q(f_reg[6]));
   DFFPOSX1 H5_reg_reg_7_ ( .CLK(clk),  .D(n1579), .Q(digest[71]));
   DFFPOSX1 f_reg_reg_7_ ( .CLK(clk),  .D(n1611), .Q(f_reg[7]));
   DFFPOSX1 H5_reg_reg_8_ ( .CLK(clk),  .D(n1578), .Q(digest[72]));
   DFFPOSX1 f_reg_reg_8_ ( .CLK(clk),  .D(n1610), .Q(f_reg[8]));
   DFFPOSX1 H5_reg_reg_9_ ( .CLK(clk),  .D(n1577), .Q(digest[73]));
   DFFPOSX1 f_reg_reg_9_ ( .CLK(clk),  .D(n1609), .Q(f_reg[9]));
   DFFPOSX1 H5_reg_reg_10_ ( .CLK(clk),  .D(n1576), .Q(digest[74]));
   DFFPOSX1 f_reg_reg_10_ ( .CLK(clk),  .D(n1608), .Q(f_reg[10]));
   DFFPOSX1 H5_reg_reg_11_ ( .CLK(clk),  .D(n1575), .Q(digest[75]));
   DFFPOSX1 f_reg_reg_11_ ( .CLK(clk),  .D(n1607), .Q(f_reg[11]));
   DFFPOSX1 H5_reg_reg_12_ ( .CLK(clk),  .D(n1574), .Q(digest[76]));
   DFFPOSX1 f_reg_reg_12_ ( .CLK(clk),  .D(n1606), .Q(f_reg[12]));
   DFFPOSX1 H5_reg_reg_13_ ( .CLK(clk),  .D(n1573), .Q(digest[77]));
   DFFPOSX1 f_reg_reg_13_ ( .CLK(clk),  .D(n1605), .Q(f_reg[13]));
   DFFPOSX1 H5_reg_reg_14_ ( .CLK(clk),  .D(n1572), .Q(digest[78]));
   DFFPOSX1 f_reg_reg_14_ ( .CLK(clk),  .D(n1604), .Q(f_reg[14]));
   DFFPOSX1 H5_reg_reg_15_ ( .CLK(clk),  .D(n1571), .Q(digest[79]));
   DFFPOSX1 f_reg_reg_15_ ( .CLK(clk),  .D(n1603), .Q(f_reg[15]));
   DFFPOSX1 H5_reg_reg_16_ ( .CLK(clk),  .D(n1570), .Q(digest[80]));
   DFFPOSX1 f_reg_reg_16_ ( .CLK(clk),  .D(n1602), .Q(f_reg[16]));
   DFFPOSX1 H5_reg_reg_17_ ( .CLK(clk),  .D(n1569), .Q(digest[81]));
   DFFPOSX1 f_reg_reg_17_ ( .CLK(clk),  .D(n1601), .Q(f_reg[17]));
   DFFPOSX1 H5_reg_reg_18_ ( .CLK(clk),  .D(n1568), .Q(digest[82]));
   DFFPOSX1 f_reg_reg_18_ ( .CLK(clk),  .D(n1600), .Q(f_reg[18]));
   DFFPOSX1 H5_reg_reg_19_ ( .CLK(clk),  .D(n1567), .Q(digest[83]));
   DFFPOSX1 f_reg_reg_19_ ( .CLK(clk),  .D(n1599), .Q(f_reg[19]));
   DFFPOSX1 H5_reg_reg_20_ ( .CLK(clk),  .D(n1566), .Q(digest[84]));
   DFFPOSX1 f_reg_reg_20_ ( .CLK(clk),  .D(n1598), .Q(f_reg[20]));
   DFFPOSX1 H5_reg_reg_21_ ( .CLK(clk),  .D(n1565), .Q(digest[85]));
   DFFPOSX1 f_reg_reg_21_ ( .CLK(clk),  .D(n1597), .Q(f_reg[21]));
   DFFPOSX1 H5_reg_reg_22_ ( .CLK(clk),  .D(n1564), .Q(digest[86]));
   DFFPOSX1 f_reg_reg_22_ ( .CLK(clk),  .D(n1596), .Q(f_reg[22]));
   DFFPOSX1 H5_reg_reg_23_ ( .CLK(clk),  .D(n1563), .Q(digest[87]));
   DFFPOSX1 f_reg_reg_23_ ( .CLK(clk),  .D(n1595), .Q(f_reg[23]));
   DFFPOSX1 H5_reg_reg_24_ ( .CLK(clk),  .D(n1562), .Q(digest[88]));
   DFFPOSX1 f_reg_reg_24_ ( .CLK(clk),  .D(n1594), .Q(f_reg[24]));
   DFFPOSX1 H5_reg_reg_25_ ( .CLK(clk),  .D(n1561), .Q(digest[89]));
   DFFPOSX1 f_reg_reg_25_ ( .CLK(clk),  .D(n1593), .Q(f_reg[25]));
   DFFPOSX1 H5_reg_reg_26_ ( .CLK(clk),  .D(n1560), .Q(digest[90]));
   DFFPOSX1 f_reg_reg_26_ ( .CLK(clk),  .D(n1592), .Q(f_reg[26]));
   DFFPOSX1 H5_reg_reg_27_ ( .CLK(clk),  .D(n1559), .Q(digest[91]));
   DFFPOSX1 f_reg_reg_27_ ( .CLK(clk),  .D(n1591), .Q(f_reg[27]));
   DFFPOSX1 H5_reg_reg_28_ ( .CLK(clk),  .D(n1558), .Q(digest[92]));
   DFFPOSX1 f_reg_reg_28_ ( .CLK(clk),  .D(n1590), .Q(f_reg[28]));
   DFFPOSX1 H5_reg_reg_29_ ( .CLK(clk),  .D(n1557), .Q(digest[93]));
   DFFPOSX1 f_reg_reg_29_ ( .CLK(clk),  .D(n1589), .Q(f_reg[29]));
   DFFPOSX1 H5_reg_reg_30_ ( .CLK(clk),  .D(n1556), .Q(digest[94]));
   DFFPOSX1 f_reg_reg_30_ ( .CLK(clk),  .D(n1588), .Q(f_reg[30]));
   DFFPOSX1 H5_reg_reg_31_ ( .CLK(clk),  .D(n1555), .Q(digest[95]));
   DFFPOSX1 g_reg_reg_31_ ( .CLK(clk),  .D(n1523), .Q(g_reg[31]));
   DFFPOSX1 H6_reg_reg_0_ ( .CLK(clk),  .D(n1522), .Q(digest[32]));
   DFFPOSX1 g_reg_reg_0_ ( .CLK(clk),  .D(n1554), .Q(g_reg[0]));
   DFFPOSX1 H6_reg_reg_1_ ( .CLK(clk),  .D(n1521), .Q(digest[33]));
   DFFPOSX1 g_reg_reg_1_ ( .CLK(clk),  .D(n1553), .Q(g_reg[1]));
   DFFPOSX1 H6_reg_reg_2_ ( .CLK(clk),  .D(n1520), .Q(digest[34]));
   DFFPOSX1 g_reg_reg_2_ ( .CLK(clk),  .D(n1552), .Q(g_reg[2]));
   DFFPOSX1 H6_reg_reg_3_ ( .CLK(clk),  .D(n1519), .Q(digest[35]));
   DFFPOSX1 g_reg_reg_3_ ( .CLK(clk),  .D(n1551), .Q(g_reg[3]));
   DFFPOSX1 H6_reg_reg_4_ ( .CLK(clk),  .D(n1518), .Q(digest[36]));
   DFFPOSX1 g_reg_reg_4_ ( .CLK(clk),  .D(n1550), .Q(g_reg[4]));
   DFFPOSX1 H6_reg_reg_5_ ( .CLK(clk),  .D(n1517), .Q(digest[37]));
   DFFPOSX1 g_reg_reg_5_ ( .CLK(clk),  .D(n1549), .Q(g_reg[5]));
   DFFPOSX1 H6_reg_reg_6_ ( .CLK(clk),  .D(n1516), .Q(digest[38]));
   DFFPOSX1 g_reg_reg_6_ ( .CLK(clk),  .D(n1548), .Q(g_reg[6]));
   DFFPOSX1 H6_reg_reg_7_ ( .CLK(clk),  .D(n1515), .Q(digest[39]));
   DFFPOSX1 g_reg_reg_7_ ( .CLK(clk),  .D(n1547), .Q(g_reg[7]));
   DFFPOSX1 H6_reg_reg_8_ ( .CLK(clk),  .D(n1514), .Q(digest[40]));
   DFFPOSX1 g_reg_reg_8_ ( .CLK(clk),  .D(n1546), .Q(g_reg[8]));
   DFFPOSX1 H6_reg_reg_9_ ( .CLK(clk),  .D(n1513), .Q(digest[41]));
   DFFPOSX1 g_reg_reg_9_ ( .CLK(clk),  .D(n1545), .Q(g_reg[9]));
   DFFPOSX1 H6_reg_reg_10_ ( .CLK(clk),  .D(n1512), .Q(digest[42]));
   DFFPOSX1 g_reg_reg_10_ ( .CLK(clk),  .D(n1544), .Q(g_reg[10]));
   DFFPOSX1 H6_reg_reg_11_ ( .CLK(clk),  .D(n1511), .Q(digest[43]));
   DFFPOSX1 g_reg_reg_11_ ( .CLK(clk),  .D(n1543), .Q(g_reg[11]));
   DFFPOSX1 H6_reg_reg_12_ ( .CLK(clk),  .D(n1510), .Q(digest[44]));
   DFFPOSX1 g_reg_reg_12_ ( .CLK(clk),  .D(n1542), .Q(g_reg[12]));
   DFFPOSX1 H6_reg_reg_13_ ( .CLK(clk),  .D(n1509), .Q(digest[45]));
   DFFPOSX1 g_reg_reg_13_ ( .CLK(clk),  .D(n1541), .Q(g_reg[13]));
   DFFPOSX1 H6_reg_reg_14_ ( .CLK(clk),  .D(n1508), .Q(digest[46]));
   DFFPOSX1 g_reg_reg_14_ ( .CLK(clk),  .D(n1540), .Q(g_reg[14]));
   DFFPOSX1 H6_reg_reg_15_ ( .CLK(clk),  .D(n1507), .Q(digest[47]));
   DFFPOSX1 g_reg_reg_15_ ( .CLK(clk),  .D(n1539), .Q(g_reg[15]));
   DFFPOSX1 H6_reg_reg_16_ ( .CLK(clk),  .D(n1506), .Q(digest[48]));
   DFFPOSX1 g_reg_reg_16_ ( .CLK(clk),  .D(n1538), .Q(g_reg[16]));
   DFFPOSX1 H6_reg_reg_17_ ( .CLK(clk),  .D(n1505), .Q(digest[49]));
   DFFPOSX1 g_reg_reg_17_ ( .CLK(clk),  .D(n1537), .Q(g_reg[17]));
   DFFPOSX1 H6_reg_reg_18_ ( .CLK(clk),  .D(n1504), .Q(digest[50]));
   DFFPOSX1 g_reg_reg_18_ ( .CLK(clk),  .D(n1536), .Q(g_reg[18]));
   DFFPOSX1 H6_reg_reg_19_ ( .CLK(clk),  .D(n1503), .Q(digest[51]));
   DFFPOSX1 g_reg_reg_19_ ( .CLK(clk),  .D(n1535), .Q(g_reg[19]));
   DFFPOSX1 H6_reg_reg_20_ ( .CLK(clk),  .D(n1502), .Q(digest[52]));
   DFFPOSX1 g_reg_reg_20_ ( .CLK(clk),  .D(n1534), .Q(g_reg[20]));
   DFFPOSX1 H6_reg_reg_21_ ( .CLK(clk),  .D(n1501), .Q(digest[53]));
   DFFPOSX1 g_reg_reg_21_ ( .CLK(clk),  .D(n1533), .Q(g_reg[21]));
   DFFPOSX1 H6_reg_reg_22_ ( .CLK(clk),  .D(n1500), .Q(digest[54]));
   DFFPOSX1 g_reg_reg_22_ ( .CLK(clk),  .D(n1532), .Q(g_reg[22]));
   DFFPOSX1 H6_reg_reg_23_ ( .CLK(clk),  .D(n1499), .Q(digest[55]));
   DFFPOSX1 g_reg_reg_23_ ( .CLK(clk),  .D(n1531), .Q(g_reg[23]));
   DFFPOSX1 H6_reg_reg_24_ ( .CLK(clk),  .D(n1498), .Q(digest[56]));
   DFFPOSX1 g_reg_reg_24_ ( .CLK(clk),  .D(n1530), .Q(g_reg[24]));
   DFFPOSX1 H6_reg_reg_25_ ( .CLK(clk),  .D(n1497), .Q(digest[57]));
   DFFPOSX1 g_reg_reg_25_ ( .CLK(clk),  .D(n1529), .Q(g_reg[25]));
   DFFPOSX1 H6_reg_reg_26_ ( .CLK(clk),  .D(n1496), .Q(digest[58]));
   DFFPOSX1 g_reg_reg_26_ ( .CLK(clk),  .D(n1528), .Q(g_reg[26]));
   DFFPOSX1 H6_reg_reg_27_ ( .CLK(clk),  .D(n1495), .Q(digest[59]));
   DFFPOSX1 g_reg_reg_27_ ( .CLK(clk),  .D(n1527), .Q(g_reg[27]));
   DFFPOSX1 H6_reg_reg_28_ ( .CLK(clk),  .D(n1494), .Q(digest[60]));
   DFFPOSX1 g_reg_reg_28_ ( .CLK(clk),  .D(n1526), .Q(g_reg[28]));
   DFFPOSX1 H6_reg_reg_29_ ( .CLK(clk),  .D(n1493), .Q(digest[61]));
   DFFPOSX1 g_reg_reg_29_ ( .CLK(clk),  .D(n1525), .Q(g_reg[29]));
   DFFPOSX1 H6_reg_reg_30_ ( .CLK(clk),  .D(n1492), .Q(digest[62]));
   DFFPOSX1 g_reg_reg_30_ ( .CLK(clk),  .D(n1524), .Q(g_reg[30]));
   DFFPOSX1 H6_reg_reg_31_ ( .CLK(clk),  .D(n1491), .Q(digest[63]));
   DFFPOSX1 h_reg_reg_31_ ( .CLK(clk),  .D(n1459), .Q(h_reg[31]));
   DFFPOSX1 H7_reg_reg_0_ ( .CLK(clk),  .D(n1458), .Q(digest[0]));
   DFFPOSX1 h_reg_reg_0_ ( .CLK(clk),  .D(n1490), .Q(h_reg[0]));
   DFFPOSX1 H7_reg_reg_1_ ( .CLK(clk),  .D(n1457), .Q(digest[1]));
   DFFPOSX1 h_reg_reg_1_ ( .CLK(clk),  .D(n1489), .Q(h_reg[1]));
   DFFPOSX1 H7_reg_reg_2_ ( .CLK(clk),  .D(n1456), .Q(digest[2]));
   DFFPOSX1 h_reg_reg_2_ ( .CLK(clk),  .D(n1488), .Q(h_reg[2]));
   DFFPOSX1 H7_reg_reg_3_ ( .CLK(clk),  .D(n1455), .Q(digest[3]));
   DFFPOSX1 h_reg_reg_3_ ( .CLK(clk),  .D(n1487), .Q(h_reg[3]));
   DFFPOSX1 H7_reg_reg_4_ ( .CLK(clk),  .D(n1454), .Q(digest[4]));
   DFFPOSX1 h_reg_reg_4_ ( .CLK(clk),  .D(n1486), .Q(h_reg[4]));
   DFFPOSX1 H7_reg_reg_5_ ( .CLK(clk),  .D(n1453), .Q(digest[5]));
   DFFPOSX1 h_reg_reg_5_ ( .CLK(clk),  .D(n1485), .Q(h_reg[5]));
   DFFPOSX1 H7_reg_reg_6_ ( .CLK(clk),  .D(n1452), .Q(digest[6]));
   DFFPOSX1 h_reg_reg_6_ ( .CLK(clk),  .D(n1484), .Q(h_reg[6]));
   DFFPOSX1 H7_reg_reg_7_ ( .CLK(clk),  .D(n1451), .Q(digest[7]));
   DFFPOSX1 h_reg_reg_7_ ( .CLK(clk),  .D(n1483), .Q(h_reg[7]));
   DFFPOSX1 H7_reg_reg_8_ ( .CLK(clk),  .D(n1450), .Q(digest[8]));
   DFFPOSX1 h_reg_reg_8_ ( .CLK(clk),  .D(n1482), .Q(h_reg[8]));
   DFFPOSX1 H7_reg_reg_9_ ( .CLK(clk),  .D(n1449), .Q(digest[9]));
   DFFPOSX1 h_reg_reg_9_ ( .CLK(clk),  .D(n1481), .Q(h_reg[9]));
   DFFPOSX1 H7_reg_reg_10_ ( .CLK(clk),  .D(n1448), .Q(digest[10]));
   DFFPOSX1 h_reg_reg_10_ ( .CLK(clk),  .D(n1480), .Q(h_reg[10]));
   DFFPOSX1 H7_reg_reg_11_ ( .CLK(clk),  .D(n1447), .Q(digest[11]));
   DFFPOSX1 h_reg_reg_11_ ( .CLK(clk),  .D(n1479), .Q(h_reg[11]));
   DFFPOSX1 H7_reg_reg_12_ ( .CLK(clk),  .D(n1446), .Q(digest[12]));
   DFFPOSX1 h_reg_reg_12_ ( .CLK(clk),  .D(n1478), .Q(h_reg[12]));
   DFFPOSX1 H7_reg_reg_13_ ( .CLK(clk),  .D(n1445), .Q(digest[13]));
   DFFPOSX1 h_reg_reg_13_ ( .CLK(clk),  .D(n1477), .Q(h_reg[13]));
   DFFPOSX1 H7_reg_reg_14_ ( .CLK(clk),  .D(n1444), .Q(digest[14]));
   DFFPOSX1 h_reg_reg_14_ ( .CLK(clk),  .D(n1476), .Q(h_reg[14]));
   DFFPOSX1 H7_reg_reg_15_ ( .CLK(clk),  .D(n1443), .Q(digest[15]));
   DFFPOSX1 h_reg_reg_15_ ( .CLK(clk),  .D(n1475), .Q(h_reg[15]));
   DFFPOSX1 H7_reg_reg_16_ ( .CLK(clk),  .D(n1442), .Q(digest[16]));
   DFFPOSX1 h_reg_reg_16_ ( .CLK(clk),  .D(n1474), .Q(h_reg[16]));
   DFFPOSX1 H7_reg_reg_17_ ( .CLK(clk),  .D(n1441), .Q(digest[17]));
   DFFPOSX1 h_reg_reg_17_ ( .CLK(clk),  .D(n1473), .Q(h_reg[17]));
   DFFPOSX1 H7_reg_reg_18_ ( .CLK(clk),  .D(n1440), .Q(digest[18]));
   DFFPOSX1 h_reg_reg_18_ ( .CLK(clk),  .D(n1472), .Q(h_reg[18]));
   DFFPOSX1 H7_reg_reg_19_ ( .CLK(clk),  .D(n1439), .Q(digest[19]));
   DFFPOSX1 h_reg_reg_19_ ( .CLK(clk),  .D(n1471), .Q(h_reg[19]));
   DFFPOSX1 H7_reg_reg_20_ ( .CLK(clk),  .D(n1438), .Q(digest[20]));
   DFFPOSX1 h_reg_reg_20_ ( .CLK(clk),  .D(n1470), .Q(h_reg[20]));
   DFFPOSX1 H7_reg_reg_21_ ( .CLK(clk),  .D(n1437), .Q(digest[21]));
   DFFPOSX1 h_reg_reg_21_ ( .CLK(clk),  .D(n1469), .Q(h_reg[21]));
   DFFPOSX1 H7_reg_reg_22_ ( .CLK(clk),  .D(n1436), .Q(digest[22]));
   DFFPOSX1 h_reg_reg_22_ ( .CLK(clk),  .D(n1468), .Q(h_reg[22]));
   DFFPOSX1 H7_reg_reg_23_ ( .CLK(clk),  .D(n1435), .Q(digest[23]));
   DFFPOSX1 h_reg_reg_23_ ( .CLK(clk),  .D(n1467), .Q(h_reg[23]));
   DFFPOSX1 H7_reg_reg_24_ ( .CLK(clk),  .D(n1434), .Q(digest[24]));
   DFFPOSX1 h_reg_reg_24_ ( .CLK(clk),  .D(n1466), .Q(h_reg[24]));
   DFFPOSX1 H7_reg_reg_25_ ( .CLK(clk),  .D(n1433), .Q(digest[25]));
   DFFPOSX1 h_reg_reg_25_ ( .CLK(clk),  .D(n1465), .Q(h_reg[25]));
   DFFPOSX1 H7_reg_reg_26_ ( .CLK(clk),  .D(n1432), .Q(digest[26]));
   DFFPOSX1 h_reg_reg_26_ ( .CLK(clk),  .D(n1464), .Q(h_reg[26]));
   DFFPOSX1 H7_reg_reg_27_ ( .CLK(clk),  .D(n1431), .Q(digest[27]));
   DFFPOSX1 h_reg_reg_27_ ( .CLK(clk),  .D(n1463), .Q(h_reg[27]));
   DFFPOSX1 H7_reg_reg_28_ ( .CLK(clk),  .D(n1430), .Q(digest[28]));
   DFFPOSX1 h_reg_reg_28_ ( .CLK(clk),  .D(n1462), .Q(h_reg[28]));
   DFFPOSX1 H7_reg_reg_29_ ( .CLK(clk),  .D(n1429), .Q(digest[29]));
   DFFPOSX1 h_reg_reg_29_ ( .CLK(clk),  .D(n1461), .Q(h_reg[29]));
   DFFPOSX1 H7_reg_reg_30_ ( .CLK(clk),  .D(n1428), .Q(digest[30]));
   DFFPOSX1 h_reg_reg_30_ ( .CLK(clk),  .D(n1460), .Q(h_reg[30]));
   DFFPOSX1 H7_reg_reg_31_ ( .CLK(clk),  .D(n1427), .Q(digest[31]));
   DFFPOSX1 a_reg_reg_31_ ( .CLK(clk),  .D(n1395), .Q(a_reg[31]));
   DFFPOSX1 H0_reg_reg_0_ ( .CLK(clk),  .D(n1394), .Q(digest[224]));
   DFFPOSX1 a_reg_reg_0_ ( .CLK(clk),  .D(n1426), .Q(a_reg[0]));
   DFFPOSX1 H0_reg_reg_1_ ( .CLK(clk),  .D(n1393), .Q(digest[225]));
   DFFPOSX1 a_reg_reg_1_ ( .CLK(clk),  .D(n1425), .Q(a_reg[1]));
   DFFPOSX1 H0_reg_reg_2_ ( .CLK(clk),  .D(n1392), .Q(digest[226]));
   DFFPOSX1 a_reg_reg_2_ ( .CLK(clk),  .D(n1424), .Q(a_reg[2]));
   DFFPOSX1 H0_reg_reg_3_ ( .CLK(clk),  .D(n1391), .Q(digest[227]));
   DFFPOSX1 a_reg_reg_3_ ( .CLK(clk),  .D(n1423), .Q(a_reg[3]));
   DFFPOSX1 H0_reg_reg_4_ ( .CLK(clk),  .D(n1390), .Q(digest[228]));
   DFFPOSX1 a_reg_reg_4_ ( .CLK(clk),  .D(n1422), .Q(a_reg[4]));
   DFFPOSX1 H0_reg_reg_5_ ( .CLK(clk),  .D(n1389), .Q(digest[229]));
   DFFPOSX1 a_reg_reg_5_ ( .CLK(clk),  .D(n1421), .Q(a_reg[5]));
   DFFPOSX1 H0_reg_reg_6_ ( .CLK(clk),  .D(n1388), .Q(digest[230]));
   DFFPOSX1 a_reg_reg_6_ ( .CLK(clk),  .D(n1420), .Q(a_reg[6]));
   DFFPOSX1 H0_reg_reg_7_ ( .CLK(clk),  .D(n1387), .Q(digest[231]));
   DFFPOSX1 a_reg_reg_7_ ( .CLK(clk),  .D(n1419), .Q(a_reg[7]));
   DFFPOSX1 H0_reg_reg_8_ ( .CLK(clk),  .D(n1386), .Q(digest[232]));
   DFFPOSX1 a_reg_reg_8_ ( .CLK(clk),  .D(n1418), .Q(a_reg[8]));
   DFFPOSX1 H0_reg_reg_9_ ( .CLK(clk),  .D(n1385), .Q(digest[233]));
   DFFPOSX1 a_reg_reg_9_ ( .CLK(clk),  .D(n1417), .Q(a_reg[9]));
   DFFPOSX1 H0_reg_reg_10_ ( .CLK(clk),  .D(n1384), .Q(digest[234]));
   DFFPOSX1 a_reg_reg_10_ ( .CLK(clk),  .D(n1416), .Q(a_reg[10]));
   DFFPOSX1 H0_reg_reg_11_ ( .CLK(clk),  .D(n1383), .Q(digest[235]));
   DFFPOSX1 a_reg_reg_11_ ( .CLK(clk),  .D(n1415), .Q(a_reg[11]));
   DFFPOSX1 H0_reg_reg_12_ ( .CLK(clk),  .D(n1382), .Q(digest[236]));
   DFFPOSX1 a_reg_reg_12_ ( .CLK(clk),  .D(n1414), .Q(a_reg[12]));
   DFFPOSX1 H0_reg_reg_13_ ( .CLK(clk),  .D(n1381), .Q(digest[237]));
   DFFPOSX1 a_reg_reg_13_ ( .CLK(clk),  .D(n1413), .Q(a_reg[13]));
   DFFPOSX1 H0_reg_reg_14_ ( .CLK(clk),  .D(n1380), .Q(digest[238]));
   DFFPOSX1 a_reg_reg_14_ ( .CLK(clk),  .D(n1412), .Q(a_reg[14]));
   DFFPOSX1 H0_reg_reg_15_ ( .CLK(clk),  .D(n1379), .Q(digest[239]));
   DFFPOSX1 a_reg_reg_15_ ( .CLK(clk),  .D(n1411), .Q(a_reg[15]));
   DFFPOSX1 H0_reg_reg_16_ ( .CLK(clk),  .D(n1378), .Q(digest[240]));
   DFFPOSX1 a_reg_reg_16_ ( .CLK(clk),  .D(n1410), .Q(a_reg[16]));
   DFFPOSX1 H0_reg_reg_17_ ( .CLK(clk),  .D(n1377), .Q(digest[241]));
   DFFPOSX1 a_reg_reg_17_ ( .CLK(clk),  .D(n1409), .Q(a_reg[17]));
   DFFPOSX1 H0_reg_reg_18_ ( .CLK(clk),  .D(n1376), .Q(digest[242]));
   DFFPOSX1 a_reg_reg_18_ ( .CLK(clk),  .D(n1408), .Q(a_reg[18]));
   DFFPOSX1 H0_reg_reg_19_ ( .CLK(clk),  .D(n1375), .Q(digest[243]));
   DFFPOSX1 a_reg_reg_19_ ( .CLK(clk),  .D(n1407), .Q(a_reg[19]));
   DFFPOSX1 H0_reg_reg_20_ ( .CLK(clk),  .D(n1374), .Q(digest[244]));
   DFFPOSX1 a_reg_reg_20_ ( .CLK(clk),  .D(n1406), .Q(a_reg[20]));
   DFFPOSX1 H0_reg_reg_21_ ( .CLK(clk),  .D(n1373), .Q(digest[245]));
   DFFPOSX1 a_reg_reg_21_ ( .CLK(clk),  .D(n1405), .Q(a_reg[21]));
   DFFPOSX1 H0_reg_reg_22_ ( .CLK(clk),  .D(n1372), .Q(digest[246]));
   DFFPOSX1 a_reg_reg_22_ ( .CLK(clk),  .D(n1404), .Q(a_reg[22]));
   DFFPOSX1 H0_reg_reg_23_ ( .CLK(clk),  .D(n1371), .Q(digest[247]));
   DFFPOSX1 a_reg_reg_23_ ( .CLK(clk),  .D(n1403), .Q(a_reg[23]));
   DFFPOSX1 H0_reg_reg_24_ ( .CLK(clk),  .D(n1370), .Q(digest[248]));
   DFFPOSX1 a_reg_reg_24_ ( .CLK(clk),  .D(n1402), .Q(a_reg[24]));
   DFFPOSX1 H0_reg_reg_25_ ( .CLK(clk),  .D(n1369), .Q(digest[249]));
   DFFPOSX1 a_reg_reg_25_ ( .CLK(clk),  .D(n1401), .Q(a_reg[25]));
   DFFPOSX1 H0_reg_reg_26_ ( .CLK(clk),  .D(n1368), .Q(digest[250]));
   DFFPOSX1 a_reg_reg_26_ ( .CLK(clk),  .D(n1400), .Q(a_reg[26]));
   DFFPOSX1 H0_reg_reg_27_ ( .CLK(clk),  .D(n1367), .Q(digest[251]));
   DFFPOSX1 a_reg_reg_27_ ( .CLK(clk),  .D(n1399), .Q(a_reg[27]));
   DFFPOSX1 H0_reg_reg_28_ ( .CLK(clk),  .D(n1366), .Q(digest[252]));
   DFFPOSX1 a_reg_reg_28_ ( .CLK(clk),  .D(n1398), .Q(a_reg[28]));
   DFFPOSX1 H0_reg_reg_29_ ( .CLK(clk),  .D(n1365), .Q(digest[253]));
   DFFPOSX1 a_reg_reg_29_ ( .CLK(clk),  .D(n1397), .Q(a_reg[29]));
   DFFPOSX1 H0_reg_reg_30_ ( .CLK(clk),  .D(n1364), .Q(digest[254]));
   DFFPOSX1 a_reg_reg_30_ ( .CLK(clk),  .D(n1396), .Q(a_reg[30]));
   DFFPOSX1 H0_reg_reg_31_ ( .CLK(clk),  .D(n1363), .Q(digest[255]));
   DFFPOSX1 b_reg_reg_31_ ( .CLK(clk),  .D(n1331), .Q(b_reg[31]));
   DFFPOSX1 H1_reg_reg_0_ ( .CLK(clk),  .D(n1330), .Q(digest[192]));
   DFFPOSX1 b_reg_reg_0_ ( .CLK(clk),  .D(n1362), .Q(b_reg[0]));
   DFFPOSX1 H1_reg_reg_1_ ( .CLK(clk),  .D(n1329), .Q(digest[193]));
   DFFPOSX1 b_reg_reg_1_ ( .CLK(clk),  .D(n1361), .Q(b_reg[1]));
   DFFPOSX1 H1_reg_reg_2_ ( .CLK(clk),  .D(n1328), .Q(digest[194]));
   DFFPOSX1 b_reg_reg_2_ ( .CLK(clk),  .D(n1360), .Q(b_reg[2]));
   DFFPOSX1 H1_reg_reg_3_ ( .CLK(clk),  .D(n1327), .Q(digest[195]));
   DFFPOSX1 b_reg_reg_3_ ( .CLK(clk),  .D(n1359), .Q(b_reg[3]));
   DFFPOSX1 H1_reg_reg_4_ ( .CLK(clk),  .D(n1326), .Q(digest[196]));
   DFFPOSX1 b_reg_reg_4_ ( .CLK(clk),  .D(n1358), .Q(b_reg[4]));
   DFFPOSX1 H1_reg_reg_5_ ( .CLK(clk),  .D(n1325), .Q(digest[197]));
   DFFPOSX1 b_reg_reg_5_ ( .CLK(clk),  .D(n1357), .Q(b_reg[5]));
   DFFPOSX1 H1_reg_reg_6_ ( .CLK(clk),  .D(n1324), .Q(digest[198]));
   DFFPOSX1 b_reg_reg_6_ ( .CLK(clk),  .D(n1356), .Q(b_reg[6]));
   DFFPOSX1 H1_reg_reg_7_ ( .CLK(clk),  .D(n1323), .Q(digest[199]));
   DFFPOSX1 b_reg_reg_7_ ( .CLK(clk),  .D(n1355), .Q(b_reg[7]));
   DFFPOSX1 H1_reg_reg_8_ ( .CLK(clk),  .D(n1322), .Q(digest[200]));
   DFFPOSX1 b_reg_reg_8_ ( .CLK(clk),  .D(n1354), .Q(b_reg[8]));
   DFFPOSX1 H1_reg_reg_9_ ( .CLK(clk),  .D(n1321), .Q(digest[201]));
   DFFPOSX1 b_reg_reg_9_ ( .CLK(clk),  .D(n1353), .Q(b_reg[9]));
   DFFPOSX1 H1_reg_reg_10_ ( .CLK(clk),  .D(n1320), .Q(digest[202]));
   DFFPOSX1 b_reg_reg_10_ ( .CLK(clk),  .D(n1352), .Q(b_reg[10]));
   DFFPOSX1 H1_reg_reg_11_ ( .CLK(clk),  .D(n1319), .Q(digest[203]));
   DFFPOSX1 b_reg_reg_11_ ( .CLK(clk),  .D(n1351), .Q(b_reg[11]));
   DFFPOSX1 H1_reg_reg_12_ ( .CLK(clk),  .D(n1318), .Q(digest[204]));
   DFFPOSX1 b_reg_reg_12_ ( .CLK(clk),  .D(n1350), .Q(b_reg[12]));
   DFFPOSX1 H1_reg_reg_13_ ( .CLK(clk),  .D(n1317), .Q(digest[205]));
   DFFPOSX1 b_reg_reg_13_ ( .CLK(clk),  .D(n1349), .Q(b_reg[13]));
   DFFPOSX1 H1_reg_reg_14_ ( .CLK(clk),  .D(n1316), .Q(digest[206]));
   DFFPOSX1 b_reg_reg_14_ ( .CLK(clk),  .D(n1348), .Q(b_reg[14]));
   DFFPOSX1 H1_reg_reg_15_ ( .CLK(clk),  .D(n1315), .Q(digest[207]));
   DFFPOSX1 b_reg_reg_15_ ( .CLK(clk),  .D(n1347), .Q(b_reg[15]));
   DFFPOSX1 H1_reg_reg_16_ ( .CLK(clk),  .D(n1314), .Q(digest[208]));
   DFFPOSX1 b_reg_reg_16_ ( .CLK(clk),  .D(n1346), .Q(b_reg[16]));
   DFFPOSX1 H1_reg_reg_17_ ( .CLK(clk),  .D(n1313), .Q(digest[209]));
   DFFPOSX1 b_reg_reg_17_ ( .CLK(clk),  .D(n1345), .Q(b_reg[17]));
   DFFPOSX1 H1_reg_reg_18_ ( .CLK(clk),  .D(n1312), .Q(digest[210]));
   DFFPOSX1 b_reg_reg_18_ ( .CLK(clk),  .D(n1344), .Q(b_reg[18]));
   DFFPOSX1 H1_reg_reg_19_ ( .CLK(clk),  .D(n1311), .Q(digest[211]));
   DFFPOSX1 b_reg_reg_19_ ( .CLK(clk),  .D(n1343), .Q(b_reg[19]));
   DFFPOSX1 H1_reg_reg_20_ ( .CLK(clk),  .D(n1310), .Q(digest[212]));
   DFFPOSX1 b_reg_reg_20_ ( .CLK(clk),  .D(n1342), .Q(b_reg[20]));
   DFFPOSX1 H1_reg_reg_21_ ( .CLK(clk),  .D(n1309), .Q(digest[213]));
   DFFPOSX1 b_reg_reg_21_ ( .CLK(clk),  .D(n1341), .Q(b_reg[21]));
   DFFPOSX1 H1_reg_reg_22_ ( .CLK(clk),  .D(n1308), .Q(digest[214]));
   DFFPOSX1 b_reg_reg_22_ ( .CLK(clk),  .D(n1340), .Q(b_reg[22]));
   DFFPOSX1 H1_reg_reg_23_ ( .CLK(clk),  .D(n1307), .Q(digest[215]));
   DFFPOSX1 b_reg_reg_23_ ( .CLK(clk),  .D(n1339), .Q(b_reg[23]));
   DFFPOSX1 H1_reg_reg_24_ ( .CLK(clk),  .D(n1306), .Q(digest[216]));
   DFFPOSX1 b_reg_reg_24_ ( .CLK(clk),  .D(n1338), .Q(b_reg[24]));
   DFFPOSX1 H1_reg_reg_25_ ( .CLK(clk),  .D(n1305), .Q(digest[217]));
   DFFPOSX1 b_reg_reg_25_ ( .CLK(clk),  .D(n1337), .Q(b_reg[25]));
   DFFPOSX1 H1_reg_reg_26_ ( .CLK(clk),  .D(n1304), .Q(digest[218]));
   DFFPOSX1 b_reg_reg_26_ ( .CLK(clk),  .D(n1336), .Q(b_reg[26]));
   DFFPOSX1 H1_reg_reg_27_ ( .CLK(clk),  .D(n1303), .Q(digest[219]));
   DFFPOSX1 b_reg_reg_27_ ( .CLK(clk),  .D(n1335), .Q(b_reg[27]));
   DFFPOSX1 H1_reg_reg_28_ ( .CLK(clk),  .D(n1302), .Q(digest[220]));
   DFFPOSX1 b_reg_reg_28_ ( .CLK(clk),  .D(n1334), .Q(b_reg[28]));
   DFFPOSX1 H1_reg_reg_29_ ( .CLK(clk),  .D(n1301), .Q(digest[221]));
   DFFPOSX1 b_reg_reg_29_ ( .CLK(clk),  .D(n1333), .Q(b_reg[29]));
   DFFPOSX1 H1_reg_reg_30_ ( .CLK(clk),  .D(n1300), .Q(digest[222]));
   DFFPOSX1 b_reg_reg_30_ ( .CLK(clk),  .D(n1332), .Q(b_reg[30]));
   DFFPOSX1 H1_reg_reg_31_ ( .CLK(clk),  .D(n1299), .Q(digest[223]));
   DFFPOSX1 c_reg_reg_31_ ( .CLK(clk),  .D(n1267), .Q(c_reg[31]));
   DFFPOSX1 H2_reg_reg_0_ ( .CLK(clk),  .D(n1266), .Q(digest[160]));
   DFFPOSX1 c_reg_reg_0_ ( .CLK(clk),  .D(n1298), .Q(c_reg[0]));
   DFFPOSX1 H2_reg_reg_1_ ( .CLK(clk),  .D(n1265), .Q(digest[161]));
   DFFPOSX1 c_reg_reg_1_ ( .CLK(clk),  .D(n1297), .Q(c_reg[1]));
   DFFPOSX1 H2_reg_reg_2_ ( .CLK(clk),  .D(n1264), .Q(digest[162]));
   DFFPOSX1 c_reg_reg_2_ ( .CLK(clk),  .D(n1296), .Q(c_reg[2]));
   DFFPOSX1 H2_reg_reg_3_ ( .CLK(clk),  .D(n1263), .Q(digest[163]));
   DFFPOSX1 c_reg_reg_3_ ( .CLK(clk),  .D(n1295), .Q(c_reg[3]));
   DFFPOSX1 H2_reg_reg_4_ ( .CLK(clk),  .D(n1262), .Q(digest[164]));
   DFFPOSX1 c_reg_reg_4_ ( .CLK(clk),  .D(n1294), .Q(c_reg[4]));
   DFFPOSX1 H2_reg_reg_5_ ( .CLK(clk),  .D(n1261), .Q(digest[165]));
   DFFPOSX1 c_reg_reg_5_ ( .CLK(clk),  .D(n1293), .Q(c_reg[5]));
   DFFPOSX1 H2_reg_reg_6_ ( .CLK(clk),  .D(n1260), .Q(digest[166]));
   DFFPOSX1 c_reg_reg_6_ ( .CLK(clk),  .D(n1292), .Q(c_reg[6]));
   DFFPOSX1 H2_reg_reg_7_ ( .CLK(clk),  .D(n1259), .Q(digest[167]));
   DFFPOSX1 c_reg_reg_7_ ( .CLK(clk),  .D(n1291), .Q(c_reg[7]));
   DFFPOSX1 H2_reg_reg_8_ ( .CLK(clk),  .D(n1258), .Q(digest[168]));
   DFFPOSX1 c_reg_reg_8_ ( .CLK(clk),  .D(n1290), .Q(c_reg[8]));
   DFFPOSX1 H2_reg_reg_9_ ( .CLK(clk),  .D(n1257), .Q(digest[169]));
   DFFPOSX1 c_reg_reg_9_ ( .CLK(clk),  .D(n1289), .Q(c_reg[9]));
   DFFPOSX1 H2_reg_reg_10_ ( .CLK(clk),  .D(n1256), .Q(digest[170]));
   DFFPOSX1 c_reg_reg_10_ ( .CLK(clk),  .D(n1288), .Q(c_reg[10]));
   DFFPOSX1 H2_reg_reg_11_ ( .CLK(clk),  .D(n1255), .Q(digest[171]));
   DFFPOSX1 c_reg_reg_11_ ( .CLK(clk),  .D(n1287), .Q(c_reg[11]));
   DFFPOSX1 H2_reg_reg_12_ ( .CLK(clk),  .D(n1254), .Q(digest[172]));
   DFFPOSX1 c_reg_reg_12_ ( .CLK(clk),  .D(n1286), .Q(c_reg[12]));
   DFFPOSX1 H2_reg_reg_13_ ( .CLK(clk),  .D(n1253), .Q(digest[173]));
   DFFPOSX1 c_reg_reg_13_ ( .CLK(clk),  .D(n1285), .Q(c_reg[13]));
   DFFPOSX1 H2_reg_reg_14_ ( .CLK(clk),  .D(n1252), .Q(digest[174]));
   DFFPOSX1 c_reg_reg_14_ ( .CLK(clk),  .D(n1284), .Q(c_reg[14]));
   DFFPOSX1 H2_reg_reg_15_ ( .CLK(clk),  .D(n1251), .Q(digest[175]));
   DFFPOSX1 c_reg_reg_15_ ( .CLK(clk),  .D(n1283), .Q(c_reg[15]));
   DFFPOSX1 H2_reg_reg_16_ ( .CLK(clk),  .D(n1250), .Q(digest[176]));
   DFFPOSX1 c_reg_reg_16_ ( .CLK(clk),  .D(n1282), .Q(c_reg[16]));
   DFFPOSX1 H2_reg_reg_17_ ( .CLK(clk),  .D(n1249), .Q(digest[177]));
   DFFPOSX1 c_reg_reg_17_ ( .CLK(clk),  .D(n1281), .Q(c_reg[17]));
   DFFPOSX1 H2_reg_reg_18_ ( .CLK(clk),  .D(n1248), .Q(digest[178]));
   DFFPOSX1 c_reg_reg_18_ ( .CLK(clk),  .D(n1280), .Q(c_reg[18]));
   DFFPOSX1 H2_reg_reg_19_ ( .CLK(clk),  .D(n1247), .Q(digest[179]));
   DFFPOSX1 c_reg_reg_19_ ( .CLK(clk),  .D(n1279), .Q(c_reg[19]));
   DFFPOSX1 H2_reg_reg_20_ ( .CLK(clk),  .D(n1246), .Q(digest[180]));
   DFFPOSX1 c_reg_reg_20_ ( .CLK(clk),  .D(n1278), .Q(c_reg[20]));
   DFFPOSX1 H2_reg_reg_21_ ( .CLK(clk),  .D(n1245), .Q(digest[181]));
   DFFPOSX1 c_reg_reg_21_ ( .CLK(clk),  .D(n1277), .Q(c_reg[21]));
   DFFPOSX1 H2_reg_reg_22_ ( .CLK(clk),  .D(n1244), .Q(digest[182]));
   DFFPOSX1 c_reg_reg_22_ ( .CLK(clk),  .D(n1276), .Q(c_reg[22]));
   DFFPOSX1 H2_reg_reg_23_ ( .CLK(clk),  .D(n1243), .Q(digest[183]));
   DFFPOSX1 c_reg_reg_23_ ( .CLK(clk),  .D(n1275), .Q(c_reg[23]));
   DFFPOSX1 H2_reg_reg_24_ ( .CLK(clk),  .D(n1242), .Q(digest[184]));
   DFFPOSX1 c_reg_reg_24_ ( .CLK(clk),  .D(n1274), .Q(c_reg[24]));
   DFFPOSX1 H2_reg_reg_25_ ( .CLK(clk),  .D(n1241), .Q(digest[185]));
   DFFPOSX1 c_reg_reg_25_ ( .CLK(clk),  .D(n1273), .Q(c_reg[25]));
   DFFPOSX1 H2_reg_reg_26_ ( .CLK(clk),  .D(n1240), .Q(digest[186]));
   DFFPOSX1 c_reg_reg_26_ ( .CLK(clk),  .D(n1272), .Q(c_reg[26]));
   DFFPOSX1 H2_reg_reg_27_ ( .CLK(clk),  .D(n1239), .Q(digest[187]));
   DFFPOSX1 c_reg_reg_27_ ( .CLK(clk),  .D(n1271), .Q(c_reg[27]));
   DFFPOSX1 H2_reg_reg_28_ ( .CLK(clk),  .D(n1238), .Q(digest[188]));
   DFFPOSX1 c_reg_reg_28_ ( .CLK(clk),  .D(n1270), .Q(c_reg[28]));
   DFFPOSX1 H2_reg_reg_29_ ( .CLK(clk),  .D(n1237), .Q(digest[189]));
   DFFPOSX1 c_reg_reg_29_ ( .CLK(clk),  .D(n1269), .Q(c_reg[29]));
   DFFPOSX1 H2_reg_reg_30_ ( .CLK(clk),  .D(n1236), .Q(digest[190]));
   DFFPOSX1 c_reg_reg_30_ ( .CLK(clk),  .D(n1268), .Q(c_reg[30]));
   DFFPOSX1 H2_reg_reg_31_ ( .CLK(clk),  .D(n1235), .Q(digest[191]));
   DFFPOSX1 d_reg_reg_31_ ( .CLK(clk),  .D(n1714), .Q(d_reg[31]));
   DFFPOSX1 H3_reg_reg_1_ ( .CLK(clk),  .D(n1713), .Q(digest[129]));
   DFFPOSX1 d_reg_reg_1_ ( .CLK(clk),  .D(n1744), .Q(d_reg[1]));
   DFFPOSX1 H3_reg_reg_2_ ( .CLK(clk),  .D(n1712), .Q(digest[130]));
   DFFPOSX1 d_reg_reg_2_ ( .CLK(clk),  .D(n1743), .Q(d_reg[2]));
   DFFPOSX1 H3_reg_reg_3_ ( .CLK(clk),  .D(n1711), .Q(digest[131]));
   DFFPOSX1 d_reg_reg_3_ ( .CLK(clk),  .D(n1742), .Q(d_reg[3]));
   DFFPOSX1 H3_reg_reg_4_ ( .CLK(clk),  .D(n1710), .Q(digest[132]));
   DFFPOSX1 d_reg_reg_4_ ( .CLK(clk),  .D(n1741), .Q(d_reg[4]));
   DFFPOSX1 H3_reg_reg_5_ ( .CLK(clk),  .D(n1709), .Q(digest[133]));
   DFFPOSX1 d_reg_reg_5_ ( .CLK(clk),  .D(n1740), .Q(d_reg[5]));
   DFFPOSX1 H3_reg_reg_6_ ( .CLK(clk),  .D(n1708), .Q(digest[134]));
   DFFPOSX1 d_reg_reg_6_ ( .CLK(clk),  .D(n1739), .Q(d_reg[6]));
   DFFPOSX1 H3_reg_reg_7_ ( .CLK(clk),  .D(n1707), .Q(digest[135]));
   DFFPOSX1 d_reg_reg_7_ ( .CLK(clk),  .D(n1738), .Q(d_reg[7]));
   DFFPOSX1 H3_reg_reg_8_ ( .CLK(clk),  .D(n1706), .Q(digest[136]));
   DFFPOSX1 d_reg_reg_8_ ( .CLK(clk),  .D(n1737), .Q(d_reg[8]));
   DFFPOSX1 H3_reg_reg_9_ ( .CLK(clk),  .D(n1705), .Q(digest[137]));
   DFFPOSX1 d_reg_reg_9_ ( .CLK(clk),  .D(n1736), .Q(d_reg[9]));
   DFFPOSX1 H3_reg_reg_10_ ( .CLK(clk),  .D(n1704), .Q(digest[138]));
   DFFPOSX1 d_reg_reg_10_ ( .CLK(clk),  .D(n1735), .Q(d_reg[10]));
   DFFPOSX1 H3_reg_reg_11_ ( .CLK(clk),  .D(n1703), .Q(digest[139]));
   DFFPOSX1 d_reg_reg_11_ ( .CLK(clk),  .D(n1734), .Q(d_reg[11]));
   DFFPOSX1 H3_reg_reg_12_ ( .CLK(clk),  .D(n1702), .Q(digest[140]));
   DFFPOSX1 d_reg_reg_12_ ( .CLK(clk),  .D(n1733), .Q(d_reg[12]));
   DFFPOSX1 H3_reg_reg_13_ ( .CLK(clk),  .D(n1701), .Q(digest[141]));
   DFFPOSX1 d_reg_reg_13_ ( .CLK(clk),  .D(n1732), .Q(d_reg[13]));
   DFFPOSX1 H3_reg_reg_14_ ( .CLK(clk),  .D(n1700), .Q(digest[142]));
   DFFPOSX1 d_reg_reg_14_ ( .CLK(clk),  .D(n1731), .Q(d_reg[14]));
   DFFPOSX1 H3_reg_reg_15_ ( .CLK(clk),  .D(n1699), .Q(digest[143]));
   DFFPOSX1 d_reg_reg_15_ ( .CLK(clk),  .D(n1730), .Q(d_reg[15]));
   DFFPOSX1 H3_reg_reg_16_ ( .CLK(clk),  .D(n1698), .Q(digest[144]));
   DFFPOSX1 d_reg_reg_16_ ( .CLK(clk),  .D(n1729), .Q(d_reg[16]));
   DFFPOSX1 H3_reg_reg_17_ ( .CLK(clk),  .D(n1697), .Q(digest[145]));
   DFFPOSX1 d_reg_reg_17_ ( .CLK(clk),  .D(n1728), .Q(d_reg[17]));
   DFFPOSX1 H3_reg_reg_18_ ( .CLK(clk),  .D(n1696), .Q(digest[146]));
   DFFPOSX1 d_reg_reg_18_ ( .CLK(clk),  .D(n1727), .Q(d_reg[18]));
   DFFPOSX1 H3_reg_reg_19_ ( .CLK(clk),  .D(n1695), .Q(digest[147]));
   DFFPOSX1 d_reg_reg_19_ ( .CLK(clk),  .D(n1726), .Q(d_reg[19]));
   DFFPOSX1 H3_reg_reg_20_ ( .CLK(clk),  .D(n1694), .Q(digest[148]));
   DFFPOSX1 d_reg_reg_20_ ( .CLK(clk),  .D(n1725), .Q(d_reg[20]));
   DFFPOSX1 H3_reg_reg_21_ ( .CLK(clk),  .D(n1693), .Q(digest[149]));
   DFFPOSX1 d_reg_reg_21_ ( .CLK(clk),  .D(n1724), .Q(d_reg[21]));
   DFFPOSX1 H3_reg_reg_22_ ( .CLK(clk),  .D(n1692), .Q(digest[150]));
   DFFPOSX1 d_reg_reg_22_ ( .CLK(clk),  .D(n1723), .Q(d_reg[22]));
   DFFPOSX1 H3_reg_reg_23_ ( .CLK(clk),  .D(n1691), .Q(digest[151]));
   DFFPOSX1 d_reg_reg_23_ ( .CLK(clk),  .D(n1722), .Q(d_reg[23]));
   DFFPOSX1 H3_reg_reg_24_ ( .CLK(clk),  .D(n1690), .Q(digest[152]));
   DFFPOSX1 d_reg_reg_24_ ( .CLK(clk),  .D(n1721), .Q(d_reg[24]));
   DFFPOSX1 H3_reg_reg_25_ ( .CLK(clk),  .D(n1689), .Q(digest[153]));
   DFFPOSX1 d_reg_reg_25_ ( .CLK(clk),  .D(n1720), .Q(d_reg[25]));
   DFFPOSX1 H3_reg_reg_26_ ( .CLK(clk),  .D(n1688), .Q(digest[154]));
   DFFPOSX1 d_reg_reg_26_ ( .CLK(clk),  .D(n1719), .Q(d_reg[26]));
   DFFPOSX1 H3_reg_reg_27_ ( .CLK(clk),  .D(n1687), .Q(digest[155]));
   DFFPOSX1 d_reg_reg_27_ ( .CLK(clk),  .D(n1718), .Q(d_reg[27]));
   DFFPOSX1 H3_reg_reg_28_ ( .CLK(clk),  .D(n1686), .Q(digest[156]));
   DFFPOSX1 d_reg_reg_28_ ( .CLK(clk),  .D(n1717), .Q(d_reg[28]));
   DFFPOSX1 H3_reg_reg_29_ ( .CLK(clk),  .D(n1685), .Q(digest[157]));
   DFFPOSX1 d_reg_reg_29_ ( .CLK(clk),  .D(n1716), .Q(d_reg[29]));
   DFFPOSX1 H3_reg_reg_30_ ( .CLK(clk),  .D(n1684), .Q(digest[158]));
   DFFPOSX1 d_reg_reg_30_ ( .CLK(clk),  .D(n1715), .Q(d_reg[30]));
   DFFPOSX1 H3_reg_reg_31_ ( .CLK(clk),  .D(n1683), .Q(digest[159]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__31_ ( .CLK(clk),  .D(w_mem_inst_n1624), .Q(w_mem_inst_w_mem[511]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__31_ ( .CLK(clk),  .D(w_mem_inst_n1656), .Q(w_mem_inst_w_mem[479]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__31_ ( .CLK(clk),  .D(w_mem_inst_n1688), .Q(w_mem_inst_w_mem[447]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__31_ ( .CLK(clk),  .D(w_mem_inst_n1720), .Q(w_mem_inst_w_mem[415]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__31_ ( .CLK(clk),  .D(w_mem_inst_n1752), .Q(w_mem_inst_w_mem[383]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__31_ ( .CLK(clk),  .D(w_mem_inst_n1784), .Q(w_mem_inst_w_mem[351]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__31_ ( .CLK(clk),  .D(w_mem_inst_n1816), .Q(w_mem_inst_w_mem[319]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__31_ ( .CLK(clk),  .D(w_mem_inst_n1848), .Q(w_mem_inst_w_mem[287]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__31_ ( .CLK(clk),  .D(w_mem_inst_n1880), .Q(w_mem_inst_w_mem[255]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__31_ ( .CLK(clk),  .D(w_mem_inst_n1912), .Q(w_mem_inst_w_mem[223]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__31_ ( .CLK(clk),  .D(w_mem_inst_n1944), .Q(w_mem_inst_w_mem[191]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__31_ ( .CLK(clk),  .D(w_mem_inst_n1976), .Q(w_mem_inst_w_mem[159]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__31_ ( .CLK(clk),  .D(w_mem_inst_n2008), .Q(w_mem_inst_w_mem[127]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__31_ ( .CLK(clk),  .D(w_mem_inst_n2040), .Q(w_mem_inst_w_mem[95]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__31_ ( .CLK(clk),  .D(w_mem_inst_n2072), .Q(w_mem_inst_w_mem[63]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__31_ ( .CLK(clk),  .D(w_mem_inst_n2104), .Q(w_mem_inst_w_mem[31]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__30_ ( .CLK(clk),  .D(w_mem_inst_n1625), .Q(w_mem_inst_w_mem[510]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__30_ ( .CLK(clk),  .D(w_mem_inst_n1657), .Q(w_mem_inst_w_mem[478]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__30_ ( .CLK(clk),  .D(w_mem_inst_n1689), .Q(w_mem_inst_w_mem[446]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__30_ ( .CLK(clk),  .D(w_mem_inst_n1721), .Q(w_mem_inst_w_mem[414]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__30_ ( .CLK(clk),  .D(w_mem_inst_n1753), .Q(w_mem_inst_w_mem[382]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__30_ ( .CLK(clk),  .D(w_mem_inst_n1785), .Q(w_mem_inst_w_mem[350]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__30_ ( .CLK(clk),  .D(w_mem_inst_n1817), .Q(w_mem_inst_w_mem[318]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__30_ ( .CLK(clk),  .D(w_mem_inst_n1849), .Q(w_mem_inst_w_mem[286]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__30_ ( .CLK(clk),  .D(w_mem_inst_n1881), .Q(w_mem_inst_w_mem[254]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__30_ ( .CLK(clk),  .D(w_mem_inst_n1913), .Q(w_mem_inst_w_mem[222]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__30_ ( .CLK(clk),  .D(w_mem_inst_n1945), .Q(w_mem_inst_w_mem[190]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__30_ ( .CLK(clk),  .D(w_mem_inst_n1977), .Q(w_mem_inst_w_mem[158]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__30_ ( .CLK(clk),  .D(w_mem_inst_n2009), .Q(w_mem_inst_w_mem[126]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__30_ ( .CLK(clk),  .D(w_mem_inst_n2041), .Q(w_mem_inst_w_mem[94]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__30_ ( .CLK(clk),  .D(w_mem_inst_n2073), .Q(w_mem_inst_w_mem[62]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__30_ ( .CLK(clk),  .D(w_mem_inst_n2105), .Q(w_mem_inst_w_mem[30]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__29_ ( .CLK(clk),  .D(w_mem_inst_n1626), .Q(w_mem_inst_w_mem[509]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__29_ ( .CLK(clk),  .D(w_mem_inst_n1658), .Q(w_mem_inst_w_mem[477]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__29_ ( .CLK(clk),  .D(w_mem_inst_n1690), .Q(w_mem_inst_w_mem[445]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__29_ ( .CLK(clk),  .D(w_mem_inst_n1722), .Q(w_mem_inst_w_mem[413]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__29_ ( .CLK(clk),  .D(w_mem_inst_n1754), .Q(w_mem_inst_w_mem[381]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__29_ ( .CLK(clk),  .D(w_mem_inst_n1786), .Q(w_mem_inst_w_mem[349]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__29_ ( .CLK(clk),  .D(w_mem_inst_n1818), .Q(w_mem_inst_w_mem[317]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__29_ ( .CLK(clk),  .D(w_mem_inst_n1850), .Q(w_mem_inst_w_mem[285]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__29_ ( .CLK(clk),  .D(w_mem_inst_n1882), .Q(w_mem_inst_w_mem[253]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__29_ ( .CLK(clk),  .D(w_mem_inst_n1914), .Q(w_mem_inst_w_mem[221]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__29_ ( .CLK(clk),  .D(w_mem_inst_n1946), .Q(w_mem_inst_w_mem[189]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__29_ ( .CLK(clk),  .D(w_mem_inst_n1978), .Q(w_mem_inst_w_mem[157]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__29_ ( .CLK(clk),  .D(w_mem_inst_n2010), .Q(w_mem_inst_w_mem[125]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__29_ ( .CLK(clk),  .D(w_mem_inst_n2042), .Q(w_mem_inst_w_mem[93]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__29_ ( .CLK(clk),  .D(w_mem_inst_n2074), .Q(w_mem_inst_w_mem[61]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__29_ ( .CLK(clk),  .D(w_mem_inst_n2106), .Q(w_mem_inst_w_mem[29]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__28_ ( .CLK(clk),  .D(w_mem_inst_n1627), .Q(w_mem_inst_w_mem[508]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__28_ ( .CLK(clk),  .D(w_mem_inst_n1659), .Q(w_mem_inst_w_mem[476]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__28_ ( .CLK(clk),  .D(w_mem_inst_n1691), .Q(w_mem_inst_w_mem[444]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__28_ ( .CLK(clk),  .D(w_mem_inst_n1723), .Q(w_mem_inst_w_mem[412]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__28_ ( .CLK(clk),  .D(w_mem_inst_n1755), .Q(w_mem_inst_w_mem[380]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__28_ ( .CLK(clk),  .D(w_mem_inst_n1787), .Q(w_mem_inst_w_mem[348]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__28_ ( .CLK(clk),  .D(w_mem_inst_n1819), .Q(w_mem_inst_w_mem[316]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__28_ ( .CLK(clk),  .D(w_mem_inst_n1851), .Q(w_mem_inst_w_mem[284]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__28_ ( .CLK(clk),  .D(w_mem_inst_n1883), .Q(w_mem_inst_w_mem[252]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__28_ ( .CLK(clk),  .D(w_mem_inst_n1915), .Q(w_mem_inst_w_mem[220]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__28_ ( .CLK(clk),  .D(w_mem_inst_n1947), .Q(w_mem_inst_w_mem[188]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__28_ ( .CLK(clk),  .D(w_mem_inst_n1979), .Q(w_mem_inst_w_mem[156]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__28_ ( .CLK(clk),  .D(w_mem_inst_n2011), .Q(w_mem_inst_w_mem[124]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__28_ ( .CLK(clk),  .D(w_mem_inst_n2043), .Q(w_mem_inst_w_mem[92]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__28_ ( .CLK(clk),  .D(w_mem_inst_n2075), .Q(w_mem_inst_w_mem[60]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__28_ ( .CLK(clk),  .D(w_mem_inst_n2107), .Q(w_mem_inst_w_mem[28]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__27_ ( .CLK(clk),  .D(w_mem_inst_n1628), .Q(w_mem_inst_w_mem[507]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__27_ ( .CLK(clk),  .D(w_mem_inst_n1660), .Q(w_mem_inst_w_mem[475]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__27_ ( .CLK(clk),  .D(w_mem_inst_n1692), .Q(w_mem_inst_w_mem[443]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__27_ ( .CLK(clk),  .D(w_mem_inst_n1724), .Q(w_mem_inst_w_mem[411]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__27_ ( .CLK(clk),  .D(w_mem_inst_n1756), .Q(w_mem_inst_w_mem[379]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__27_ ( .CLK(clk),  .D(w_mem_inst_n1788), .Q(w_mem_inst_w_mem[347]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__27_ ( .CLK(clk),  .D(w_mem_inst_n1820), .Q(w_mem_inst_w_mem[315]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__27_ ( .CLK(clk),  .D(w_mem_inst_n1852), .Q(w_mem_inst_w_mem[283]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__27_ ( .CLK(clk),  .D(w_mem_inst_n1884), .Q(w_mem_inst_w_mem[251]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__27_ ( .CLK(clk),  .D(w_mem_inst_n1916), .Q(w_mem_inst_w_mem[219]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__27_ ( .CLK(clk),  .D(w_mem_inst_n1948), .Q(w_mem_inst_w_mem[187]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__27_ ( .CLK(clk),  .D(w_mem_inst_n1980), .Q(w_mem_inst_w_mem[155]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__27_ ( .CLK(clk),  .D(w_mem_inst_n2012), .Q(w_mem_inst_w_mem[123]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__27_ ( .CLK(clk),  .D(w_mem_inst_n2044), .Q(w_mem_inst_w_mem[91]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__27_ ( .CLK(clk),  .D(w_mem_inst_n2076), .Q(w_mem_inst_w_mem[59]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__27_ ( .CLK(clk),  .D(w_mem_inst_n2108), .Q(w_mem_inst_w_mem[27]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__26_ ( .CLK(clk),  .D(w_mem_inst_n1629), .Q(w_mem_inst_w_mem[506]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__26_ ( .CLK(clk),  .D(w_mem_inst_n1661), .Q(w_mem_inst_w_mem[474]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__26_ ( .CLK(clk),  .D(w_mem_inst_n1693), .Q(w_mem_inst_w_mem[442]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__26_ ( .CLK(clk),  .D(w_mem_inst_n1725), .Q(w_mem_inst_w_mem[410]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__26_ ( .CLK(clk),  .D(w_mem_inst_n1757), .Q(w_mem_inst_w_mem[378]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__26_ ( .CLK(clk),  .D(w_mem_inst_n1789), .Q(w_mem_inst_w_mem[346]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__26_ ( .CLK(clk),  .D(w_mem_inst_n1821), .Q(w_mem_inst_w_mem[314]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__26_ ( .CLK(clk),  .D(w_mem_inst_n1853), .Q(w_mem_inst_w_mem[282]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__26_ ( .CLK(clk),  .D(w_mem_inst_n1885), .Q(w_mem_inst_w_mem[250]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__26_ ( .CLK(clk),  .D(w_mem_inst_n1917), .Q(w_mem_inst_w_mem[218]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__26_ ( .CLK(clk),  .D(w_mem_inst_n1949), .Q(w_mem_inst_w_mem[186]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__26_ ( .CLK(clk),  .D(w_mem_inst_n1981), .Q(w_mem_inst_w_mem[154]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__26_ ( .CLK(clk),  .D(w_mem_inst_n2013), .Q(w_mem_inst_w_mem[122]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__26_ ( .CLK(clk),  .D(w_mem_inst_n2045), .Q(w_mem_inst_w_mem[90]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__26_ ( .CLK(clk),  .D(w_mem_inst_n2077), .Q(w_mem_inst_w_mem[58]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__26_ ( .CLK(clk),  .D(w_mem_inst_n2109), .Q(w_mem_inst_w_mem[26]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__25_ ( .CLK(clk),  .D(w_mem_inst_n1630), .Q(w_mem_inst_w_mem[505]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__25_ ( .CLK(clk),  .D(w_mem_inst_n1662), .Q(w_mem_inst_w_mem[473]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__25_ ( .CLK(clk),  .D(w_mem_inst_n1694), .Q(w_mem_inst_w_mem[441]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__25_ ( .CLK(clk),  .D(w_mem_inst_n1726), .Q(w_mem_inst_w_mem[409]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__25_ ( .CLK(clk),  .D(w_mem_inst_n1758), .Q(w_mem_inst_w_mem[377]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__25_ ( .CLK(clk),  .D(w_mem_inst_n1790), .Q(w_mem_inst_w_mem[345]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__25_ ( .CLK(clk),  .D(w_mem_inst_n1822), .Q(w_mem_inst_w_mem[313]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__25_ ( .CLK(clk),  .D(w_mem_inst_n1854), .Q(w_mem_inst_w_mem[281]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__25_ ( .CLK(clk),  .D(w_mem_inst_n1886), .Q(w_mem_inst_w_mem[249]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__25_ ( .CLK(clk),  .D(w_mem_inst_n1918), .Q(w_mem_inst_w_mem[217]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__25_ ( .CLK(clk),  .D(w_mem_inst_n1950), .Q(w_mem_inst_w_mem[185]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__25_ ( .CLK(clk),  .D(w_mem_inst_n1982), .Q(w_mem_inst_w_mem[153]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__25_ ( .CLK(clk),  .D(w_mem_inst_n2014), .Q(w_mem_inst_w_mem[121]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__25_ ( .CLK(clk),  .D(w_mem_inst_n2046), .Q(w_mem_inst_w_mem[89]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__25_ ( .CLK(clk),  .D(w_mem_inst_n2078), .Q(w_mem_inst_w_mem[57]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__25_ ( .CLK(clk),  .D(w_mem_inst_n2110), .Q(w_mem_inst_w_mem[25]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__24_ ( .CLK(clk),  .D(w_mem_inst_n1631), .Q(w_mem_inst_w_mem[504]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__24_ ( .CLK(clk),  .D(w_mem_inst_n1663), .Q(w_mem_inst_w_mem[472]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__24_ ( .CLK(clk),  .D(w_mem_inst_n1695), .Q(w_mem_inst_w_mem[440]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__24_ ( .CLK(clk),  .D(w_mem_inst_n1727), .Q(w_mem_inst_w_mem[408]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__24_ ( .CLK(clk),  .D(w_mem_inst_n1759), .Q(w_mem_inst_w_mem[376]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__24_ ( .CLK(clk),  .D(w_mem_inst_n1791), .Q(w_mem_inst_w_mem[344]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__24_ ( .CLK(clk),  .D(w_mem_inst_n1823), .Q(w_mem_inst_w_mem[312]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__24_ ( .CLK(clk),  .D(w_mem_inst_n1855), .Q(w_mem_inst_w_mem[280]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__24_ ( .CLK(clk),  .D(w_mem_inst_n1887), .Q(w_mem_inst_w_mem[248]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__24_ ( .CLK(clk),  .D(w_mem_inst_n1919), .Q(w_mem_inst_w_mem[216]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__24_ ( .CLK(clk),  .D(w_mem_inst_n1951), .Q(w_mem_inst_w_mem[184]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__24_ ( .CLK(clk),  .D(w_mem_inst_n1983), .Q(w_mem_inst_w_mem[152]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__24_ ( .CLK(clk),  .D(w_mem_inst_n2015), .Q(w_mem_inst_w_mem[120]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__24_ ( .CLK(clk),  .D(w_mem_inst_n2047), .Q(w_mem_inst_w_mem[88]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__24_ ( .CLK(clk),  .D(w_mem_inst_n2079), .Q(w_mem_inst_w_mem[56]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__24_ ( .CLK(clk),  .D(w_mem_inst_n2111), .Q(w_mem_inst_w_mem[24]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__23_ ( .CLK(clk),  .D(w_mem_inst_n1632), .Q(w_mem_inst_w_mem[503]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__23_ ( .CLK(clk),  .D(w_mem_inst_n1664), .Q(w_mem_inst_w_mem[471]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__23_ ( .CLK(clk),  .D(w_mem_inst_n1696), .Q(w_mem_inst_w_mem[439]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__23_ ( .CLK(clk),  .D(w_mem_inst_n1728), .Q(w_mem_inst_w_mem[407]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__23_ ( .CLK(clk),  .D(w_mem_inst_n1760), .Q(w_mem_inst_w_mem[375]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__23_ ( .CLK(clk),  .D(w_mem_inst_n1792), .Q(w_mem_inst_w_mem[343]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__23_ ( .CLK(clk),  .D(w_mem_inst_n1824), .Q(w_mem_inst_w_mem[311]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__23_ ( .CLK(clk),  .D(w_mem_inst_n1856), .Q(w_mem_inst_w_mem[279]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__23_ ( .CLK(clk),  .D(w_mem_inst_n1888), .Q(w_mem_inst_w_mem[247]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__23_ ( .CLK(clk),  .D(w_mem_inst_n1920), .Q(w_mem_inst_w_mem[215]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__23_ ( .CLK(clk),  .D(w_mem_inst_n1952), .Q(w_mem_inst_w_mem[183]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__23_ ( .CLK(clk),  .D(w_mem_inst_n1984), .Q(w_mem_inst_w_mem[151]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__23_ ( .CLK(clk),  .D(w_mem_inst_n2016), .Q(w_mem_inst_w_mem[119]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__23_ ( .CLK(clk),  .D(w_mem_inst_n2048), .Q(w_mem_inst_w_mem[87]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__23_ ( .CLK(clk),  .D(w_mem_inst_n2080), .Q(w_mem_inst_w_mem[55]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__23_ ( .CLK(clk),  .D(w_mem_inst_n2112), .Q(w_mem_inst_w_mem[23]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__22_ ( .CLK(clk),  .D(w_mem_inst_n1633), .Q(w_mem_inst_w_mem[502]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__22_ ( .CLK(clk),  .D(w_mem_inst_n1665), .Q(w_mem_inst_w_mem[470]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__22_ ( .CLK(clk),  .D(w_mem_inst_n1697), .Q(w_mem_inst_w_mem[438]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__22_ ( .CLK(clk),  .D(w_mem_inst_n1729), .Q(w_mem_inst_w_mem[406]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__22_ ( .CLK(clk),  .D(w_mem_inst_n1761), .Q(w_mem_inst_w_mem[374]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__22_ ( .CLK(clk),  .D(w_mem_inst_n1793), .Q(w_mem_inst_w_mem[342]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__22_ ( .CLK(clk),  .D(w_mem_inst_n1825), .Q(w_mem_inst_w_mem[310]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__22_ ( .CLK(clk),  .D(w_mem_inst_n1857), .Q(w_mem_inst_w_mem[278]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__22_ ( .CLK(clk),  .D(w_mem_inst_n1889), .Q(w_mem_inst_w_mem[246]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__22_ ( .CLK(clk),  .D(w_mem_inst_n1921), .Q(w_mem_inst_w_mem[214]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__22_ ( .CLK(clk),  .D(w_mem_inst_n1953), .Q(w_mem_inst_w_mem[182]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__22_ ( .CLK(clk),  .D(w_mem_inst_n1985), .Q(w_mem_inst_w_mem[150]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__22_ ( .CLK(clk),  .D(w_mem_inst_n2017), .Q(w_mem_inst_w_mem[118]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__22_ ( .CLK(clk),  .D(w_mem_inst_n2049), .Q(w_mem_inst_w_mem[86]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__22_ ( .CLK(clk),  .D(w_mem_inst_n2081), .Q(w_mem_inst_w_mem[54]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__22_ ( .CLK(clk),  .D(w_mem_inst_n2113), .Q(w_mem_inst_w_mem[22]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__21_ ( .CLK(clk),  .D(w_mem_inst_n1634), .Q(w_mem_inst_w_mem[501]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__21_ ( .CLK(clk),  .D(w_mem_inst_n1666), .Q(w_mem_inst_w_mem[469]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__21_ ( .CLK(clk),  .D(w_mem_inst_n1698), .Q(w_mem_inst_w_mem[437]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__21_ ( .CLK(clk),  .D(w_mem_inst_n1730), .Q(w_mem_inst_w_mem[405]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__21_ ( .CLK(clk),  .D(w_mem_inst_n1762), .Q(w_mem_inst_w_mem[373]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__21_ ( .CLK(clk),  .D(w_mem_inst_n1794), .Q(w_mem_inst_w_mem[341]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__21_ ( .CLK(clk),  .D(w_mem_inst_n1826), .Q(w_mem_inst_w_mem[309]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__21_ ( .CLK(clk),  .D(w_mem_inst_n1858), .Q(w_mem_inst_w_mem[277]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__21_ ( .CLK(clk),  .D(w_mem_inst_n1890), .Q(w_mem_inst_w_mem[245]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__21_ ( .CLK(clk),  .D(w_mem_inst_n1922), .Q(w_mem_inst_w_mem[213]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__21_ ( .CLK(clk),  .D(w_mem_inst_n1954), .Q(w_mem_inst_w_mem[181]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__21_ ( .CLK(clk),  .D(w_mem_inst_n1986), .Q(w_mem_inst_w_mem[149]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__21_ ( .CLK(clk),  .D(w_mem_inst_n2018), .Q(w_mem_inst_w_mem[117]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__21_ ( .CLK(clk),  .D(w_mem_inst_n2050), .Q(w_mem_inst_w_mem[85]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__21_ ( .CLK(clk),  .D(w_mem_inst_n2082), .Q(w_mem_inst_w_mem[53]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__21_ ( .CLK(clk),  .D(w_mem_inst_n2114), .Q(w_mem_inst_w_mem[21]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__20_ ( .CLK(clk),  .D(w_mem_inst_n1635), .Q(w_mem_inst_w_mem[500]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__20_ ( .CLK(clk),  .D(w_mem_inst_n1667), .Q(w_mem_inst_w_mem[468]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__20_ ( .CLK(clk),  .D(w_mem_inst_n1699), .Q(w_mem_inst_w_mem[436]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__20_ ( .CLK(clk),  .D(w_mem_inst_n1731), .Q(w_mem_inst_w_mem[404]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__20_ ( .CLK(clk),  .D(w_mem_inst_n1763), .Q(w_mem_inst_w_mem[372]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__20_ ( .CLK(clk),  .D(w_mem_inst_n1795), .Q(w_mem_inst_w_mem[340]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__20_ ( .CLK(clk),  .D(w_mem_inst_n1827), .Q(w_mem_inst_w_mem[308]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__20_ ( .CLK(clk),  .D(w_mem_inst_n1859), .Q(w_mem_inst_w_mem[276]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__20_ ( .CLK(clk),  .D(w_mem_inst_n1891), .Q(w_mem_inst_w_mem[244]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__20_ ( .CLK(clk),  .D(w_mem_inst_n1923), .Q(w_mem_inst_w_mem[212]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__20_ ( .CLK(clk),  .D(w_mem_inst_n1955), .Q(w_mem_inst_w_mem[180]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__20_ ( .CLK(clk),  .D(w_mem_inst_n1987), .Q(w_mem_inst_w_mem[148]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__20_ ( .CLK(clk),  .D(w_mem_inst_n2019), .Q(w_mem_inst_w_mem[116]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__20_ ( .CLK(clk),  .D(w_mem_inst_n2051), .Q(w_mem_inst_w_mem[84]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__20_ ( .CLK(clk),  .D(w_mem_inst_n2083), .Q(w_mem_inst_w_mem[52]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__20_ ( .CLK(clk),  .D(w_mem_inst_n2115), .Q(w_mem_inst_w_mem[20]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__19_ ( .CLK(clk),  .D(w_mem_inst_n1636), .Q(w_mem_inst_w_mem[499]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__19_ ( .CLK(clk),  .D(w_mem_inst_n1668), .Q(w_mem_inst_w_mem[467]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__19_ ( .CLK(clk),  .D(w_mem_inst_n1700), .Q(w_mem_inst_w_mem[435]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__19_ ( .CLK(clk),  .D(w_mem_inst_n1732), .Q(w_mem_inst_w_mem[403]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__19_ ( .CLK(clk),  .D(w_mem_inst_n1764), .Q(w_mem_inst_w_mem[371]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__19_ ( .CLK(clk),  .D(w_mem_inst_n1796), .Q(w_mem_inst_w_mem[339]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__19_ ( .CLK(clk),  .D(w_mem_inst_n1828), .Q(w_mem_inst_w_mem[307]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__19_ ( .CLK(clk),  .D(w_mem_inst_n1860), .Q(w_mem_inst_w_mem[275]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__19_ ( .CLK(clk),  .D(w_mem_inst_n1892), .Q(w_mem_inst_w_mem[243]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__19_ ( .CLK(clk),  .D(w_mem_inst_n1924), .Q(w_mem_inst_w_mem[211]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__19_ ( .CLK(clk),  .D(w_mem_inst_n1956), .Q(w_mem_inst_w_mem[179]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__19_ ( .CLK(clk),  .D(w_mem_inst_n1988), .Q(w_mem_inst_w_mem[147]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__19_ ( .CLK(clk),  .D(w_mem_inst_n2020), .Q(w_mem_inst_w_mem[115]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__19_ ( .CLK(clk),  .D(w_mem_inst_n2052), .Q(w_mem_inst_w_mem[83]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__19_ ( .CLK(clk),  .D(w_mem_inst_n2084), .Q(w_mem_inst_w_mem[51]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__19_ ( .CLK(clk),  .D(w_mem_inst_n2116), .Q(w_mem_inst_w_mem[19]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__18_ ( .CLK(clk),  .D(w_mem_inst_n1637), .Q(w_mem_inst_w_mem[498]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__18_ ( .CLK(clk),  .D(w_mem_inst_n1669), .Q(w_mem_inst_w_mem[466]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__18_ ( .CLK(clk),  .D(w_mem_inst_n1701), .Q(w_mem_inst_w_mem[434]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__18_ ( .CLK(clk),  .D(w_mem_inst_n1733), .Q(w_mem_inst_w_mem[402]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__18_ ( .CLK(clk),  .D(w_mem_inst_n1765), .Q(w_mem_inst_w_mem[370]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__18_ ( .CLK(clk),  .D(w_mem_inst_n1797), .Q(w_mem_inst_w_mem[338]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__18_ ( .CLK(clk),  .D(w_mem_inst_n1829), .Q(w_mem_inst_w_mem[306]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__18_ ( .CLK(clk),  .D(w_mem_inst_n1861), .Q(w_mem_inst_w_mem[274]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__18_ ( .CLK(clk),  .D(w_mem_inst_n1893), .Q(w_mem_inst_w_mem[242]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__18_ ( .CLK(clk),  .D(w_mem_inst_n1925), .Q(w_mem_inst_w_mem[210]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__18_ ( .CLK(clk),  .D(w_mem_inst_n1957), .Q(w_mem_inst_w_mem[178]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__18_ ( .CLK(clk),  .D(w_mem_inst_n1989), .Q(w_mem_inst_w_mem[146]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__18_ ( .CLK(clk),  .D(w_mem_inst_n2021), .Q(w_mem_inst_w_mem[114]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__18_ ( .CLK(clk),  .D(w_mem_inst_n2053), .Q(w_mem_inst_w_mem[82]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__18_ ( .CLK(clk),  .D(w_mem_inst_n2085), .Q(w_mem_inst_w_mem[50]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__18_ ( .CLK(clk),  .D(w_mem_inst_n2117), .Q(w_mem_inst_w_mem[18]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__17_ ( .CLK(clk),  .D(w_mem_inst_n1638), .Q(w_mem_inst_w_mem[497]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__17_ ( .CLK(clk),  .D(w_mem_inst_n1670), .Q(w_mem_inst_w_mem[465]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__17_ ( .CLK(clk),  .D(w_mem_inst_n1702), .Q(w_mem_inst_w_mem[433]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__17_ ( .CLK(clk),  .D(w_mem_inst_n1734), .Q(w_mem_inst_w_mem[401]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__17_ ( .CLK(clk),  .D(w_mem_inst_n1766), .Q(w_mem_inst_w_mem[369]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__17_ ( .CLK(clk),  .D(w_mem_inst_n1798), .Q(w_mem_inst_w_mem[337]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__17_ ( .CLK(clk),  .D(w_mem_inst_n1830), .Q(w_mem_inst_w_mem[305]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__17_ ( .CLK(clk),  .D(w_mem_inst_n1862), .Q(w_mem_inst_w_mem[273]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__17_ ( .CLK(clk),  .D(w_mem_inst_n1894), .Q(w_mem_inst_w_mem[241]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__17_ ( .CLK(clk),  .D(w_mem_inst_n1926), .Q(w_mem_inst_w_mem[209]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__17_ ( .CLK(clk),  .D(w_mem_inst_n1958), .Q(w_mem_inst_w_mem[177]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__17_ ( .CLK(clk),  .D(w_mem_inst_n1990), .Q(w_mem_inst_w_mem[145]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__17_ ( .CLK(clk),  .D(w_mem_inst_n2022), .Q(w_mem_inst_w_mem[113]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__17_ ( .CLK(clk),  .D(w_mem_inst_n2054), .Q(w_mem_inst_w_mem[81]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__17_ ( .CLK(clk),  .D(w_mem_inst_n2086), .Q(w_mem_inst_w_mem[49]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__17_ ( .CLK(clk),  .D(w_mem_inst_n2118), .Q(w_mem_inst_w_mem[17]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__16_ ( .CLK(clk),  .D(w_mem_inst_n1639), .Q(w_mem_inst_w_mem[496]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__16_ ( .CLK(clk),  .D(w_mem_inst_n1671), .Q(w_mem_inst_w_mem[464]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__16_ ( .CLK(clk),  .D(w_mem_inst_n1703), .Q(w_mem_inst_w_mem[432]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__16_ ( .CLK(clk),  .D(w_mem_inst_n1735), .Q(w_mem_inst_w_mem[400]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__16_ ( .CLK(clk),  .D(w_mem_inst_n1767), .Q(w_mem_inst_w_mem[368]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__16_ ( .CLK(clk),  .D(w_mem_inst_n1799), .Q(w_mem_inst_w_mem[336]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__16_ ( .CLK(clk),  .D(w_mem_inst_n1831), .Q(w_mem_inst_w_mem[304]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__16_ ( .CLK(clk),  .D(w_mem_inst_n1863), .Q(w_mem_inst_w_mem[272]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__16_ ( .CLK(clk),  .D(w_mem_inst_n1895), .Q(w_mem_inst_w_mem[240]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__16_ ( .CLK(clk),  .D(w_mem_inst_n1927), .Q(w_mem_inst_w_mem[208]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__16_ ( .CLK(clk),  .D(w_mem_inst_n1959), .Q(w_mem_inst_w_mem[176]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__16_ ( .CLK(clk),  .D(w_mem_inst_n1991), .Q(w_mem_inst_w_mem[144]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__16_ ( .CLK(clk),  .D(w_mem_inst_n2023), .Q(w_mem_inst_w_mem[112]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__16_ ( .CLK(clk),  .D(w_mem_inst_n2055), .Q(w_mem_inst_w_mem[80]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__16_ ( .CLK(clk),  .D(w_mem_inst_n2087), .Q(w_mem_inst_w_mem[48]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__16_ ( .CLK(clk),  .D(w_mem_inst_n2119), .Q(w_mem_inst_w_mem[16]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__15_ ( .CLK(clk),  .D(w_mem_inst_n1640), .Q(w_mem_inst_w_mem[495]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__15_ ( .CLK(clk),  .D(w_mem_inst_n1672), .Q(w_mem_inst_w_mem[463]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__15_ ( .CLK(clk),  .D(w_mem_inst_n1704), .Q(w_mem_inst_w_mem[431]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__15_ ( .CLK(clk),  .D(w_mem_inst_n1736), .Q(w_mem_inst_w_mem[399]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__15_ ( .CLK(clk),  .D(w_mem_inst_n1768), .Q(w_mem_inst_w_mem[367]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__15_ ( .CLK(clk),  .D(w_mem_inst_n1800), .Q(w_mem_inst_w_mem[335]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__15_ ( .CLK(clk),  .D(w_mem_inst_n1832), .Q(w_mem_inst_w_mem[303]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__15_ ( .CLK(clk),  .D(w_mem_inst_n1864), .Q(w_mem_inst_w_mem[271]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__15_ ( .CLK(clk),  .D(w_mem_inst_n1896), .Q(w_mem_inst_w_mem[239]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__15_ ( .CLK(clk),  .D(w_mem_inst_n1928), .Q(w_mem_inst_w_mem[207]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__15_ ( .CLK(clk),  .D(w_mem_inst_n1960), .Q(w_mem_inst_w_mem[175]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__15_ ( .CLK(clk),  .D(w_mem_inst_n1992), .Q(w_mem_inst_w_mem[143]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__15_ ( .CLK(clk),  .D(w_mem_inst_n2024), .Q(w_mem_inst_w_mem[111]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__15_ ( .CLK(clk),  .D(w_mem_inst_n2056), .Q(w_mem_inst_w_mem[79]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__15_ ( .CLK(clk),  .D(w_mem_inst_n2088), .Q(w_mem_inst_w_mem[47]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__15_ ( .CLK(clk),  .D(w_mem_inst_n2120), .Q(w_mem_inst_w_mem[15]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__14_ ( .CLK(clk),  .D(w_mem_inst_n1641), .Q(w_mem_inst_w_mem[494]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__14_ ( .CLK(clk),  .D(w_mem_inst_n1673), .Q(w_mem_inst_w_mem[462]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__14_ ( .CLK(clk),  .D(w_mem_inst_n1705), .Q(w_mem_inst_w_mem[430]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__14_ ( .CLK(clk),  .D(w_mem_inst_n1737), .Q(w_mem_inst_w_mem[398]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__14_ ( .CLK(clk),  .D(w_mem_inst_n1769), .Q(w_mem_inst_w_mem[366]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__14_ ( .CLK(clk),  .D(w_mem_inst_n1801), .Q(w_mem_inst_w_mem[334]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__14_ ( .CLK(clk),  .D(w_mem_inst_n1833), .Q(w_mem_inst_w_mem[302]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__14_ ( .CLK(clk),  .D(w_mem_inst_n1865), .Q(w_mem_inst_w_mem[270]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__14_ ( .CLK(clk),  .D(w_mem_inst_n1897), .Q(w_mem_inst_w_mem[238]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__14_ ( .CLK(clk),  .D(w_mem_inst_n1929), .Q(w_mem_inst_w_mem[206]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__14_ ( .CLK(clk),  .D(w_mem_inst_n1961), .Q(w_mem_inst_w_mem[174]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__14_ ( .CLK(clk),  .D(w_mem_inst_n1993), .Q(w_mem_inst_w_mem[142]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__14_ ( .CLK(clk),  .D(w_mem_inst_n2025), .Q(w_mem_inst_w_mem[110]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__14_ ( .CLK(clk),  .D(w_mem_inst_n2057), .Q(w_mem_inst_w_mem[78]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__14_ ( .CLK(clk),  .D(w_mem_inst_n2089), .Q(w_mem_inst_w_mem[46]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__14_ ( .CLK(clk),  .D(w_mem_inst_n2121), .Q(w_mem_inst_w_mem[14]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__13_ ( .CLK(clk),  .D(w_mem_inst_n1642), .Q(w_mem_inst_w_mem[493]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__13_ ( .CLK(clk),  .D(w_mem_inst_n1674), .Q(w_mem_inst_w_mem[461]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__13_ ( .CLK(clk),  .D(w_mem_inst_n1706), .Q(w_mem_inst_w_mem[429]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__13_ ( .CLK(clk),  .D(w_mem_inst_n1738), .Q(w_mem_inst_w_mem[397]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__13_ ( .CLK(clk),  .D(w_mem_inst_n1770), .Q(w_mem_inst_w_mem[365]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__13_ ( .CLK(clk),  .D(w_mem_inst_n1802), .Q(w_mem_inst_w_mem[333]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__13_ ( .CLK(clk),  .D(w_mem_inst_n1834), .Q(w_mem_inst_w_mem[301]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__13_ ( .CLK(clk),  .D(w_mem_inst_n1866), .Q(w_mem_inst_w_mem[269]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__13_ ( .CLK(clk),  .D(w_mem_inst_n1898), .Q(w_mem_inst_w_mem[237]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__13_ ( .CLK(clk),  .D(w_mem_inst_n1930), .Q(w_mem_inst_w_mem[205]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__13_ ( .CLK(clk),  .D(w_mem_inst_n1962), .Q(w_mem_inst_w_mem[173]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__13_ ( .CLK(clk),  .D(w_mem_inst_n1994), .Q(w_mem_inst_w_mem[141]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__13_ ( .CLK(clk),  .D(w_mem_inst_n2026), .Q(w_mem_inst_w_mem[109]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__13_ ( .CLK(clk),  .D(w_mem_inst_n2058), .Q(w_mem_inst_w_mem[77]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__13_ ( .CLK(clk),  .D(w_mem_inst_n2090), .Q(w_mem_inst_w_mem[45]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__13_ ( .CLK(clk),  .D(w_mem_inst_n2122), .Q(w_mem_inst_w_mem[13]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__12_ ( .CLK(clk),  .D(w_mem_inst_n1643), .Q(w_mem_inst_w_mem[492]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__12_ ( .CLK(clk),  .D(w_mem_inst_n1675), .Q(w_mem_inst_w_mem[460]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__12_ ( .CLK(clk),  .D(w_mem_inst_n1707), .Q(w_mem_inst_w_mem[428]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__12_ ( .CLK(clk),  .D(w_mem_inst_n1739), .Q(w_mem_inst_w_mem[396]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__12_ ( .CLK(clk),  .D(w_mem_inst_n1771), .Q(w_mem_inst_w_mem[364]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__12_ ( .CLK(clk),  .D(w_mem_inst_n1803), .Q(w_mem_inst_w_mem[332]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__12_ ( .CLK(clk),  .D(w_mem_inst_n1835), .Q(w_mem_inst_w_mem[300]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__12_ ( .CLK(clk),  .D(w_mem_inst_n1867), .Q(w_mem_inst_w_mem[268]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__12_ ( .CLK(clk),  .D(w_mem_inst_n1899), .Q(w_mem_inst_w_mem[236]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__12_ ( .CLK(clk),  .D(w_mem_inst_n1931), .Q(w_mem_inst_w_mem[204]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__12_ ( .CLK(clk),  .D(w_mem_inst_n1963), .Q(w_mem_inst_w_mem[172]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__12_ ( .CLK(clk),  .D(w_mem_inst_n1995), .Q(w_mem_inst_w_mem[140]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__12_ ( .CLK(clk),  .D(w_mem_inst_n2027), .Q(w_mem_inst_w_mem[108]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__12_ ( .CLK(clk),  .D(w_mem_inst_n2059), .Q(w_mem_inst_w_mem[76]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__12_ ( .CLK(clk),  .D(w_mem_inst_n2091), .Q(w_mem_inst_w_mem[44]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__12_ ( .CLK(clk),  .D(w_mem_inst_n2123), .Q(w_mem_inst_w_mem[12]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__11_ ( .CLK(clk),  .D(w_mem_inst_n1644), .Q(w_mem_inst_w_mem[491]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__11_ ( .CLK(clk),  .D(w_mem_inst_n1676), .Q(w_mem_inst_w_mem[459]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__11_ ( .CLK(clk),  .D(w_mem_inst_n1708), .Q(w_mem_inst_w_mem[427]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__11_ ( .CLK(clk),  .D(w_mem_inst_n1740), .Q(w_mem_inst_w_mem[395]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__11_ ( .CLK(clk),  .D(w_mem_inst_n1772), .Q(w_mem_inst_w_mem[363]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__11_ ( .CLK(clk),  .D(w_mem_inst_n1804), .Q(w_mem_inst_w_mem[331]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__11_ ( .CLK(clk),  .D(w_mem_inst_n1836), .Q(w_mem_inst_w_mem[299]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__11_ ( .CLK(clk),  .D(w_mem_inst_n1868), .Q(w_mem_inst_w_mem[267]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__11_ ( .CLK(clk),  .D(w_mem_inst_n1900), .Q(w_mem_inst_w_mem[235]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__11_ ( .CLK(clk),  .D(w_mem_inst_n1932), .Q(w_mem_inst_w_mem[203]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__11_ ( .CLK(clk),  .D(w_mem_inst_n1964), .Q(w_mem_inst_w_mem[171]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__11_ ( .CLK(clk),  .D(w_mem_inst_n1996), .Q(w_mem_inst_w_mem[139]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__11_ ( .CLK(clk),  .D(w_mem_inst_n2028), .Q(w_mem_inst_w_mem[107]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__11_ ( .CLK(clk),  .D(w_mem_inst_n2060), .Q(w_mem_inst_w_mem[75]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__11_ ( .CLK(clk),  .D(w_mem_inst_n2092), .Q(w_mem_inst_w_mem[43]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__11_ ( .CLK(clk),  .D(w_mem_inst_n2124), .Q(w_mem_inst_w_mem[11]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__10_ ( .CLK(clk),  .D(w_mem_inst_n1645), .Q(w_mem_inst_w_mem[490]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__10_ ( .CLK(clk),  .D(w_mem_inst_n1677), .Q(w_mem_inst_w_mem[458]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__10_ ( .CLK(clk),  .D(w_mem_inst_n1709), .Q(w_mem_inst_w_mem[426]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__10_ ( .CLK(clk),  .D(w_mem_inst_n1741), .Q(w_mem_inst_w_mem[394]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__10_ ( .CLK(clk),  .D(w_mem_inst_n1773), .Q(w_mem_inst_w_mem[362]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__10_ ( .CLK(clk),  .D(w_mem_inst_n1805), .Q(w_mem_inst_w_mem[330]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__10_ ( .CLK(clk),  .D(w_mem_inst_n1837), .Q(w_mem_inst_w_mem[298]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__10_ ( .CLK(clk),  .D(w_mem_inst_n1869), .Q(w_mem_inst_w_mem[266]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__10_ ( .CLK(clk),  .D(w_mem_inst_n1901), .Q(w_mem_inst_w_mem[234]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__10_ ( .CLK(clk),  .D(w_mem_inst_n1933), .Q(w_mem_inst_w_mem[202]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__10_ ( .CLK(clk),  .D(w_mem_inst_n1965), .Q(w_mem_inst_w_mem[170]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__10_ ( .CLK(clk),  .D(w_mem_inst_n1997), .Q(w_mem_inst_w_mem[138]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__10_ ( .CLK(clk),  .D(w_mem_inst_n2029), .Q(w_mem_inst_w_mem[106]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__10_ ( .CLK(clk),  .D(w_mem_inst_n2061), .Q(w_mem_inst_w_mem[74]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__10_ ( .CLK(clk),  .D(w_mem_inst_n2093), .Q(w_mem_inst_w_mem[42]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__10_ ( .CLK(clk),  .D(w_mem_inst_n2125), .Q(w_mem_inst_w_mem[10]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__9_ ( .CLK(clk),  .D(w_mem_inst_n1646), .Q(w_mem_inst_w_mem[489]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__9_ ( .CLK(clk),  .D(w_mem_inst_n1678), .Q(w_mem_inst_w_mem[457]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__9_ ( .CLK(clk),  .D(w_mem_inst_n1710), .Q(w_mem_inst_w_mem[425]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__9_ ( .CLK(clk),  .D(w_mem_inst_n1742), .Q(w_mem_inst_w_mem[393]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__9_ ( .CLK(clk),  .D(w_mem_inst_n1774), .Q(w_mem_inst_w_mem[361]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__9_ ( .CLK(clk),  .D(w_mem_inst_n1806), .Q(w_mem_inst_w_mem[329]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__9_ ( .CLK(clk),  .D(w_mem_inst_n1838), .Q(w_mem_inst_w_mem[297]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__9_ ( .CLK(clk),  .D(w_mem_inst_n1870), .Q(w_mem_inst_w_mem[265]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__9_ ( .CLK(clk),  .D(w_mem_inst_n1902), .Q(w_mem_inst_w_mem[233]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__9_ ( .CLK(clk),  .D(w_mem_inst_n1934), .Q(w_mem_inst_w_mem[201]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__9_ ( .CLK(clk),  .D(w_mem_inst_n1966), .Q(w_mem_inst_w_mem[169]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__9_ ( .CLK(clk),  .D(w_mem_inst_n1998), .Q(w_mem_inst_w_mem[137]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__9_ ( .CLK(clk),  .D(w_mem_inst_n2030), .Q(w_mem_inst_w_mem[105]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__9_ ( .CLK(clk),  .D(w_mem_inst_n2062), .Q(w_mem_inst_w_mem[73]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__9_ ( .CLK(clk),  .D(w_mem_inst_n2094), .Q(w_mem_inst_w_mem[41]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__9_ ( .CLK(clk),  .D(w_mem_inst_n2126), .Q(w_mem_inst_w_mem[9]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__8_ ( .CLK(clk),  .D(w_mem_inst_n1647), .Q(w_mem_inst_w_mem[488]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__8_ ( .CLK(clk),  .D(w_mem_inst_n1679), .Q(w_mem_inst_w_mem[456]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__8_ ( .CLK(clk),  .D(w_mem_inst_n1711), .Q(w_mem_inst_w_mem[424]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__8_ ( .CLK(clk),  .D(w_mem_inst_n1743), .Q(w_mem_inst_w_mem[392]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__8_ ( .CLK(clk),  .D(w_mem_inst_n1775), .Q(w_mem_inst_w_mem[360]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__8_ ( .CLK(clk),  .D(w_mem_inst_n1807), .Q(w_mem_inst_w_mem[328]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__8_ ( .CLK(clk),  .D(w_mem_inst_n1839), .Q(w_mem_inst_w_mem[296]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__8_ ( .CLK(clk),  .D(w_mem_inst_n1871), .Q(w_mem_inst_w_mem[264]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__8_ ( .CLK(clk),  .D(w_mem_inst_n1903), .Q(w_mem_inst_w_mem[232]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__8_ ( .CLK(clk),  .D(w_mem_inst_n1935), .Q(w_mem_inst_w_mem[200]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__8_ ( .CLK(clk),  .D(w_mem_inst_n1967), .Q(w_mem_inst_w_mem[168]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__8_ ( .CLK(clk),  .D(w_mem_inst_n1999), .Q(w_mem_inst_w_mem[136]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__8_ ( .CLK(clk),  .D(w_mem_inst_n2031), .Q(w_mem_inst_w_mem[104]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__8_ ( .CLK(clk),  .D(w_mem_inst_n2063), .Q(w_mem_inst_w_mem[72]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__8_ ( .CLK(clk),  .D(w_mem_inst_n2095), .Q(w_mem_inst_w_mem[40]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__8_ ( .CLK(clk),  .D(w_mem_inst_n2127), .Q(w_mem_inst_w_mem[8]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__7_ ( .CLK(clk),  .D(w_mem_inst_n1648), .Q(w_mem_inst_w_mem[487]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__7_ ( .CLK(clk),  .D(w_mem_inst_n1680), .Q(w_mem_inst_w_mem[455]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__7_ ( .CLK(clk),  .D(w_mem_inst_n1712), .Q(w_mem_inst_w_mem[423]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__7_ ( .CLK(clk),  .D(w_mem_inst_n1744), .Q(w_mem_inst_w_mem[391]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__7_ ( .CLK(clk),  .D(w_mem_inst_n1776), .Q(w_mem_inst_w_mem[359]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__7_ ( .CLK(clk),  .D(w_mem_inst_n1808), .Q(w_mem_inst_w_mem[327]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__7_ ( .CLK(clk),  .D(w_mem_inst_n1840), .Q(w_mem_inst_w_mem[295]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__7_ ( .CLK(clk),  .D(w_mem_inst_n1872), .Q(w_mem_inst_w_mem[263]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__7_ ( .CLK(clk),  .D(w_mem_inst_n1904), .Q(w_mem_inst_w_mem[231]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__7_ ( .CLK(clk),  .D(w_mem_inst_n1936), .Q(w_mem_inst_w_mem[199]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__7_ ( .CLK(clk),  .D(w_mem_inst_n1968), .Q(w_mem_inst_w_mem[167]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__7_ ( .CLK(clk),  .D(w_mem_inst_n2000), .Q(w_mem_inst_w_mem[135]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__7_ ( .CLK(clk),  .D(w_mem_inst_n2032), .Q(w_mem_inst_w_mem[103]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__7_ ( .CLK(clk),  .D(w_mem_inst_n2064), .Q(w_mem_inst_w_mem[71]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__7_ ( .CLK(clk),  .D(w_mem_inst_n2096), .Q(w_mem_inst_w_mem[39]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__7_ ( .CLK(clk),  .D(w_mem_inst_n2128), .Q(w_mem_inst_w_mem[7]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__6_ ( .CLK(clk),  .D(w_mem_inst_n1649), .Q(w_mem_inst_w_mem[486]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__6_ ( .CLK(clk),  .D(w_mem_inst_n1681), .Q(w_mem_inst_w_mem[454]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__6_ ( .CLK(clk),  .D(w_mem_inst_n1713), .Q(w_mem_inst_w_mem[422]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__6_ ( .CLK(clk),  .D(w_mem_inst_n1745), .Q(w_mem_inst_w_mem[390]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__6_ ( .CLK(clk),  .D(w_mem_inst_n1777), .Q(w_mem_inst_w_mem[358]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__6_ ( .CLK(clk),  .D(w_mem_inst_n1809), .Q(w_mem_inst_w_mem[326]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__6_ ( .CLK(clk),  .D(w_mem_inst_n1841), .Q(w_mem_inst_w_mem[294]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__6_ ( .CLK(clk),  .D(w_mem_inst_n1873), .Q(w_mem_inst_w_mem[262]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__6_ ( .CLK(clk),  .D(w_mem_inst_n1905), .Q(w_mem_inst_w_mem[230]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__6_ ( .CLK(clk),  .D(w_mem_inst_n1937), .Q(w_mem_inst_w_mem[198]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__6_ ( .CLK(clk),  .D(w_mem_inst_n1969), .Q(w_mem_inst_w_mem[166]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__6_ ( .CLK(clk),  .D(w_mem_inst_n2001), .Q(w_mem_inst_w_mem[134]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__6_ ( .CLK(clk),  .D(w_mem_inst_n2033), .Q(w_mem_inst_w_mem[102]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__6_ ( .CLK(clk),  .D(w_mem_inst_n2065), .Q(w_mem_inst_w_mem[70]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__6_ ( .CLK(clk),  .D(w_mem_inst_n2097), .Q(w_mem_inst_w_mem[38]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__6_ ( .CLK(clk),  .D(w_mem_inst_n2129), .Q(w_mem_inst_w_mem[6]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__5_ ( .CLK(clk),  .D(w_mem_inst_n1650), .Q(w_mem_inst_w_mem[485]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__5_ ( .CLK(clk),  .D(w_mem_inst_n1682), .Q(w_mem_inst_w_mem[453]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__5_ ( .CLK(clk),  .D(w_mem_inst_n1714), .Q(w_mem_inst_w_mem[421]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__5_ ( .CLK(clk),  .D(w_mem_inst_n1746), .Q(w_mem_inst_w_mem[389]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__5_ ( .CLK(clk),  .D(w_mem_inst_n1778), .Q(w_mem_inst_w_mem[357]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__5_ ( .CLK(clk),  .D(w_mem_inst_n1810), .Q(w_mem_inst_w_mem[325]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__5_ ( .CLK(clk),  .D(w_mem_inst_n1842), .Q(w_mem_inst_w_mem[293]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__5_ ( .CLK(clk),  .D(w_mem_inst_n1874), .Q(w_mem_inst_w_mem[261]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__5_ ( .CLK(clk),  .D(w_mem_inst_n1906), .Q(w_mem_inst_w_mem[229]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__5_ ( .CLK(clk),  .D(w_mem_inst_n1938), .Q(w_mem_inst_w_mem[197]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__5_ ( .CLK(clk),  .D(w_mem_inst_n1970), .Q(w_mem_inst_w_mem[165]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__5_ ( .CLK(clk),  .D(w_mem_inst_n2002), .Q(w_mem_inst_w_mem[133]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__5_ ( .CLK(clk),  .D(w_mem_inst_n2034), .Q(w_mem_inst_w_mem[101]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__5_ ( .CLK(clk),  .D(w_mem_inst_n2066), .Q(w_mem_inst_w_mem[69]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__5_ ( .CLK(clk),  .D(w_mem_inst_n2098), .Q(w_mem_inst_w_mem[37]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__5_ ( .CLK(clk),  .D(w_mem_inst_n2130), .Q(w_mem_inst_w_mem[5]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__4_ ( .CLK(clk),  .D(w_mem_inst_n1651), .Q(w_mem_inst_w_mem[484]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__4_ ( .CLK(clk),  .D(w_mem_inst_n1683), .Q(w_mem_inst_w_mem[452]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__4_ ( .CLK(clk),  .D(w_mem_inst_n1715), .Q(w_mem_inst_w_mem[420]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__4_ ( .CLK(clk),  .D(w_mem_inst_n1747), .Q(w_mem_inst_w_mem[388]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__4_ ( .CLK(clk),  .D(w_mem_inst_n1779), .Q(w_mem_inst_w_mem[356]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__4_ ( .CLK(clk),  .D(w_mem_inst_n1811), .Q(w_mem_inst_w_mem[324]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__4_ ( .CLK(clk),  .D(w_mem_inst_n1843), .Q(w_mem_inst_w_mem[292]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__4_ ( .CLK(clk),  .D(w_mem_inst_n1875), .Q(w_mem_inst_w_mem[260]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__4_ ( .CLK(clk),  .D(w_mem_inst_n1907), .Q(w_mem_inst_w_mem[228]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__4_ ( .CLK(clk),  .D(w_mem_inst_n1939), .Q(w_mem_inst_w_mem[196]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__4_ ( .CLK(clk),  .D(w_mem_inst_n1971), .Q(w_mem_inst_w_mem[164]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__4_ ( .CLK(clk),  .D(w_mem_inst_n2003), .Q(w_mem_inst_w_mem[132]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__4_ ( .CLK(clk),  .D(w_mem_inst_n2035), .Q(w_mem_inst_w_mem[100]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__4_ ( .CLK(clk),  .D(w_mem_inst_n2067), .Q(w_mem_inst_w_mem[68]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__4_ ( .CLK(clk),  .D(w_mem_inst_n2099), .Q(w_mem_inst_w_mem[36]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__4_ ( .CLK(clk),  .D(w_mem_inst_n2131), .Q(w_mem_inst_w_mem[4]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__3_ ( .CLK(clk),  .D(w_mem_inst_n1652), .Q(w_mem_inst_w_mem[483]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__3_ ( .CLK(clk),  .D(w_mem_inst_n1684), .Q(w_mem_inst_w_mem[451]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__3_ ( .CLK(clk),  .D(w_mem_inst_n1716), .Q(w_mem_inst_w_mem[419]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__3_ ( .CLK(clk),  .D(w_mem_inst_n1748), .Q(w_mem_inst_w_mem[387]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__3_ ( .CLK(clk),  .D(w_mem_inst_n1780), .Q(w_mem_inst_w_mem[355]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__3_ ( .CLK(clk),  .D(w_mem_inst_n1812), .Q(w_mem_inst_w_mem[323]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__3_ ( .CLK(clk),  .D(w_mem_inst_n1844), .Q(w_mem_inst_w_mem[291]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__3_ ( .CLK(clk),  .D(w_mem_inst_n1876), .Q(w_mem_inst_w_mem[259]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__3_ ( .CLK(clk),  .D(w_mem_inst_n1908), .Q(w_mem_inst_w_mem[227]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__3_ ( .CLK(clk),  .D(w_mem_inst_n1940), .Q(w_mem_inst_w_mem[195]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__3_ ( .CLK(clk),  .D(w_mem_inst_n1972), .Q(w_mem_inst_w_mem[163]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__3_ ( .CLK(clk),  .D(w_mem_inst_n2004), .Q(w_mem_inst_w_mem[131]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__3_ ( .CLK(clk),  .D(w_mem_inst_n2036), .Q(w_mem_inst_w_mem[99]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__3_ ( .CLK(clk),  .D(w_mem_inst_n2068), .Q(w_mem_inst_w_mem[67]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__3_ ( .CLK(clk),  .D(w_mem_inst_n2100), .Q(w_mem_inst_w_mem[35]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__3_ ( .CLK(clk),  .D(w_mem_inst_n2132), .Q(w_mem_inst_w_mem[3]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__2_ ( .CLK(clk),  .D(w_mem_inst_n1653), .Q(w_mem_inst_w_mem[482]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__2_ ( .CLK(clk),  .D(w_mem_inst_n1685), .Q(w_mem_inst_w_mem[450]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__2_ ( .CLK(clk),  .D(w_mem_inst_n1717), .Q(w_mem_inst_w_mem[418]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__2_ ( .CLK(clk),  .D(w_mem_inst_n1749), .Q(w_mem_inst_w_mem[386]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__2_ ( .CLK(clk),  .D(w_mem_inst_n1781), .Q(w_mem_inst_w_mem[354]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__2_ ( .CLK(clk),  .D(w_mem_inst_n1813), .Q(w_mem_inst_w_mem[322]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__2_ ( .CLK(clk),  .D(w_mem_inst_n1845), .Q(w_mem_inst_w_mem[290]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__2_ ( .CLK(clk),  .D(w_mem_inst_n1877), .Q(w_mem_inst_w_mem[258]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__2_ ( .CLK(clk),  .D(w_mem_inst_n1909), .Q(w_mem_inst_w_mem[226]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__2_ ( .CLK(clk),  .D(w_mem_inst_n1941), .Q(w_mem_inst_w_mem[194]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__2_ ( .CLK(clk),  .D(w_mem_inst_n1973), .Q(w_mem_inst_w_mem[162]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__2_ ( .CLK(clk),  .D(w_mem_inst_n2005), .Q(w_mem_inst_w_mem[130]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__2_ ( .CLK(clk),  .D(w_mem_inst_n2037), .Q(w_mem_inst_w_mem[98]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__2_ ( .CLK(clk),  .D(w_mem_inst_n2069), .Q(w_mem_inst_w_mem[66]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__2_ ( .CLK(clk),  .D(w_mem_inst_n2101), .Q(w_mem_inst_w_mem[34]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__2_ ( .CLK(clk),  .D(w_mem_inst_n2133), .Q(w_mem_inst_w_mem[2]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__1_ ( .CLK(clk),  .D(w_mem_inst_n1654), .Q(w_mem_inst_w_mem[481]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__1_ ( .CLK(clk),  .D(w_mem_inst_n1686), .Q(w_mem_inst_w_mem[449]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__1_ ( .CLK(clk),  .D(w_mem_inst_n1718), .Q(w_mem_inst_w_mem[417]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__1_ ( .CLK(clk),  .D(w_mem_inst_n1750), .Q(w_mem_inst_w_mem[385]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__1_ ( .CLK(clk),  .D(w_mem_inst_n1782), .Q(w_mem_inst_w_mem[353]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__1_ ( .CLK(clk),  .D(w_mem_inst_n1814), .Q(w_mem_inst_w_mem[321]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__1_ ( .CLK(clk),  .D(w_mem_inst_n1846), .Q(w_mem_inst_w_mem[289]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__1_ ( .CLK(clk),  .D(w_mem_inst_n1878), .Q(w_mem_inst_w_mem[257]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__1_ ( .CLK(clk),  .D(w_mem_inst_n1910), .Q(w_mem_inst_w_mem[225]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__1_ ( .CLK(clk),  .D(w_mem_inst_n1942), .Q(w_mem_inst_w_mem[193]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__1_ ( .CLK(clk),  .D(w_mem_inst_n1974), .Q(w_mem_inst_w_mem[161]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__1_ ( .CLK(clk),  .D(w_mem_inst_n2006), .Q(w_mem_inst_w_mem[129]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__1_ ( .CLK(clk),  .D(w_mem_inst_n2038), .Q(w_mem_inst_w_mem[97]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__1_ ( .CLK(clk),  .D(w_mem_inst_n2070), .Q(w_mem_inst_w_mem[65]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__1_ ( .CLK(clk),  .D(w_mem_inst_n2102), .Q(w_mem_inst_w_mem[33]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__1_ ( .CLK(clk),  .D(w_mem_inst_n2134), .Q(w_mem_inst_w_mem[1]));
   DFFPOSX1 w_mem_inst_w_mem_reg_0__0_ ( .CLK(clk),  .D(w_mem_inst_n1655), .Q(w_mem_inst_w_mem[480]));
   DFFPOSX1 w_mem_inst_w_mem_reg_1__0_ ( .CLK(clk),  .D(w_mem_inst_n1687), .Q(w_mem_inst_w_mem[448]));
   DFFPOSX1 w_mem_inst_w_mem_reg_2__0_ ( .CLK(clk),  .D(w_mem_inst_n1719), .Q(w_mem_inst_w_mem[416]));
   DFFPOSX1 w_mem_inst_w_mem_reg_3__0_ ( .CLK(clk),  .D(w_mem_inst_n1751), .Q(w_mem_inst_w_mem[384]));
   DFFPOSX1 w_mem_inst_w_mem_reg_4__0_ ( .CLK(clk),  .D(w_mem_inst_n1783), .Q(w_mem_inst_w_mem[352]));
   DFFPOSX1 w_mem_inst_w_mem_reg_5__0_ ( .CLK(clk),  .D(w_mem_inst_n1815), .Q(w_mem_inst_w_mem[320]));
   DFFPOSX1 w_mem_inst_w_mem_reg_6__0_ ( .CLK(clk),  .D(w_mem_inst_n1847), .Q(w_mem_inst_w_mem[288]));
   DFFPOSX1 w_mem_inst_w_mem_reg_7__0_ ( .CLK(clk),  .D(w_mem_inst_n1879), .Q(w_mem_inst_w_mem[256]));
   DFFPOSX1 w_mem_inst_w_mem_reg_8__0_ ( .CLK(clk),  .D(w_mem_inst_n1911), .Q(w_mem_inst_w_mem[224]));
   DFFPOSX1 w_mem_inst_w_mem_reg_9__0_ ( .CLK(clk),  .D(w_mem_inst_n1943), .Q(w_mem_inst_w_mem[192]));
   DFFPOSX1 w_mem_inst_w_mem_reg_10__0_ ( .CLK(clk),  .D(w_mem_inst_n1975), .Q(w_mem_inst_w_mem[160]));
   DFFPOSX1 w_mem_inst_w_mem_reg_11__0_ ( .CLK(clk),  .D(w_mem_inst_n2007), .Q(w_mem_inst_w_mem[128]));
   DFFPOSX1 w_mem_inst_w_mem_reg_12__0_ ( .CLK(clk),  .D(w_mem_inst_n2039), .Q(w_mem_inst_w_mem[96]));
   DFFPOSX1 w_mem_inst_w_mem_reg_13__0_ ( .CLK(clk),  .D(w_mem_inst_n2071), .Q(w_mem_inst_w_mem[64]));
   DFFPOSX1 w_mem_inst_w_mem_reg_14__0_ ( .CLK(clk),  .D(w_mem_inst_n2103), .Q(w_mem_inst_w_mem[32]));
   DFFPOSX1 w_mem_inst_w_mem_reg_15__0_ ( .CLK(clk),  .D(w_mem_inst_n2135), .Q(w_mem_inst_w_mem[0]));
   DFFPOSX1 w_mem_inst_w_ctr_reg_reg_4_ ( .CLK(clk),  .D(w_mem_inst_n2136), .Q(w_mem_inst_w_ctr_reg[4]));
   DFFPOSX1 w_mem_inst_w_ctr_reg_reg_3_ ( .CLK(clk),  .D(w_mem_inst_n2137), .Q(w_mem_inst_w_ctr_reg[3]));
   DFFPOSX1 w_mem_inst_w_ctr_reg_reg_2_ ( .CLK(clk),  .D(w_mem_inst_n2138), .Q(w_mem_inst_w_ctr_reg[2]));
   DFFPOSX1 w_mem_inst_w_ctr_reg_reg_1_ ( .CLK(clk),  .D(w_mem_inst_n2139), .Q(w_mem_inst_w_ctr_reg[1]));
   DFFPOSX1 w_mem_inst_w_ctr_reg_reg_5_ ( .CLK(clk),  .D(w_mem_inst_n2141), .Q(w_mem_inst_w_ctr_reg[5]));
   DFFPOSX1 w_mem_inst_sha256_w_mem_ctrl_reg_reg_0_ ( .CLK(clk),  .D(w_mem_inst_n2140), .Q(w_mem_inst_sha256_w_mem_ctrl_reg_0_));
   DFFPOSX1 w_mem_inst_w_ctr_reg_reg_0_ ( .CLK(clk),  .D(w_mem_inst_n2142), .Q(w_mem_inst_w_ctr_reg[0]));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_1 ( .A(w_mem_inst_N638),  .B(w_mem_inst_w_mem[193]),  .C(n2964), .YC(w_mem_inst_add_2_root_add_945_3_carry[2]), .YS(w_mem_inst_N641));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_2 ( .A(w_mem_inst_N637),  .B(w_mem_inst_w_mem[194]),  .C(w_mem_inst_add_2_root_add_945_3_carry[2]), .YC(w_mem_inst_add_2_root_add_945_3_carry[3]), .YS(w_mem_inst_N642));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_3 ( .A(w_mem_inst_N636),  .B(w_mem_inst_w_mem[195]),  .C(w_mem_inst_add_2_root_add_945_3_carry[3]), .YC(w_mem_inst_add_2_root_add_945_3_carry[4]), .YS(w_mem_inst_N643));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_4 ( .A(w_mem_inst_N635),  .B(w_mem_inst_w_mem[196]),  .C(w_mem_inst_add_2_root_add_945_3_carry[4]), .YC(w_mem_inst_add_2_root_add_945_3_carry[5]), .YS(w_mem_inst_N644));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_5 ( .A(w_mem_inst_N634),  .B(w_mem_inst_w_mem[197]),  .C(w_mem_inst_add_2_root_add_945_3_carry[5]), .YC(w_mem_inst_add_2_root_add_945_3_carry[6]), .YS(w_mem_inst_N645));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_6 ( .A(w_mem_inst_N633),  .B(w_mem_inst_w_mem[198]),  .C(w_mem_inst_add_2_root_add_945_3_carry[6]), .YC(w_mem_inst_add_2_root_add_945_3_carry[7]), .YS(w_mem_inst_N646));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_7 ( .A(w_mem_inst_N632),  .B(w_mem_inst_w_mem[199]),  .C(w_mem_inst_add_2_root_add_945_3_carry[7]), .YC(w_mem_inst_add_2_root_add_945_3_carry[8]), .YS(w_mem_inst_N647));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_8 ( .A(w_mem_inst_N631),  .B(w_mem_inst_w_mem[200]),  .C(w_mem_inst_add_2_root_add_945_3_carry[8]), .YC(w_mem_inst_add_2_root_add_945_3_carry[9]), .YS(w_mem_inst_N648));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_9 ( .A(w_mem_inst_N630),  .B(w_mem_inst_w_mem[201]),  .C(w_mem_inst_add_2_root_add_945_3_carry[9]), .YC(w_mem_inst_add_2_root_add_945_3_carry[10]), .YS(w_mem_inst_N649));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_10 ( .A(w_mem_inst_N629),  .B(w_mem_inst_w_mem[202]),  .C(w_mem_inst_add_2_root_add_945_3_carry[10]), .YC(w_mem_inst_add_2_root_add_945_3_carry[11]), .YS(w_mem_inst_N650));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_11 ( .A(w_mem_inst_N628),  .B(w_mem_inst_w_mem[203]),  .C(w_mem_inst_add_2_root_add_945_3_carry[11]), .YC(w_mem_inst_add_2_root_add_945_3_carry[12]), .YS(w_mem_inst_N651));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_12 ( .A(w_mem_inst_N627),  .B(w_mem_inst_w_mem[204]),  .C(w_mem_inst_add_2_root_add_945_3_carry[12]), .YC(w_mem_inst_add_2_root_add_945_3_carry[13]), .YS(w_mem_inst_N652));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_13 ( .A(w_mem_inst_N626),  .B(w_mem_inst_w_mem[205]),  .C(w_mem_inst_add_2_root_add_945_3_carry[13]), .YC(w_mem_inst_add_2_root_add_945_3_carry[14]), .YS(w_mem_inst_N653));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_14 ( .A(w_mem_inst_N625),  .B(w_mem_inst_w_mem[206]),  .C(w_mem_inst_add_2_root_add_945_3_carry[14]), .YC(w_mem_inst_add_2_root_add_945_3_carry[15]), .YS(w_mem_inst_N654));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_15 ( .A(w_mem_inst_N624),  .B(w_mem_inst_w_mem[207]),  .C(w_mem_inst_add_2_root_add_945_3_carry[15]), .YC(w_mem_inst_add_2_root_add_945_3_carry[16]), .YS(w_mem_inst_N655));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_16 ( .A(w_mem_inst_N623),  .B(w_mem_inst_w_mem[208]),  .C(w_mem_inst_add_2_root_add_945_3_carry[16]), .YC(w_mem_inst_add_2_root_add_945_3_carry[17]), .YS(w_mem_inst_N656));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_17 ( .A(w_mem_inst_N622),  .B(w_mem_inst_w_mem[209]),  .C(w_mem_inst_add_2_root_add_945_3_carry[17]), .YC(w_mem_inst_add_2_root_add_945_3_carry[18]), .YS(w_mem_inst_N657));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_18 ( .A(w_mem_inst_N621),  .B(w_mem_inst_w_mem[210]),  .C(w_mem_inst_add_2_root_add_945_3_carry[18]), .YC(w_mem_inst_add_2_root_add_945_3_carry[19]), .YS(w_mem_inst_N658));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_19 ( .A(w_mem_inst_N620),  .B(w_mem_inst_w_mem[211]),  .C(w_mem_inst_add_2_root_add_945_3_carry[19]), .YC(w_mem_inst_add_2_root_add_945_3_carry[20]), .YS(w_mem_inst_N659));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_20 ( .A(w_mem_inst_N619),  .B(w_mem_inst_w_mem[212]),  .C(w_mem_inst_add_2_root_add_945_3_carry[20]), .YC(w_mem_inst_add_2_root_add_945_3_carry[21]), .YS(w_mem_inst_N660));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_21 ( .A(w_mem_inst_N618),  .B(w_mem_inst_w_mem[213]),  .C(w_mem_inst_add_2_root_add_945_3_carry[21]), .YC(w_mem_inst_add_2_root_add_945_3_carry[22]), .YS(w_mem_inst_N661));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_22 ( .A(w_mem_inst_N617),  .B(w_mem_inst_w_mem[214]),  .C(w_mem_inst_add_2_root_add_945_3_carry[22]), .YC(w_mem_inst_add_2_root_add_945_3_carry[23]), .YS(w_mem_inst_N662));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_23 ( .A(w_mem_inst_N616),  .B(w_mem_inst_w_mem[215]),  .C(w_mem_inst_add_2_root_add_945_3_carry[23]), .YC(w_mem_inst_add_2_root_add_945_3_carry[24]), .YS(w_mem_inst_N663));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_24 ( .A(w_mem_inst_N615),  .B(w_mem_inst_w_mem[216]),  .C(w_mem_inst_add_2_root_add_945_3_carry[24]), .YC(w_mem_inst_add_2_root_add_945_3_carry[25]), .YS(w_mem_inst_N664));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_25 ( .A(w_mem_inst_N614),  .B(w_mem_inst_w_mem[217]),  .C(w_mem_inst_add_2_root_add_945_3_carry[25]), .YC(w_mem_inst_add_2_root_add_945_3_carry[26]), .YS(w_mem_inst_N665));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_26 ( .A(w_mem_inst_N613),  .B(w_mem_inst_w_mem[218]),  .C(w_mem_inst_add_2_root_add_945_3_carry[26]), .YC(w_mem_inst_add_2_root_add_945_3_carry[27]), .YS(w_mem_inst_N666));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_27 ( .A(w_mem_inst_N612),  .B(w_mem_inst_w_mem[219]),  .C(w_mem_inst_add_2_root_add_945_3_carry[27]), .YC(w_mem_inst_add_2_root_add_945_3_carry[28]), .YS(w_mem_inst_N667));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_28 ( .A(w_mem_inst_N611),  .B(w_mem_inst_w_mem[220]),  .C(w_mem_inst_add_2_root_add_945_3_carry[28]), .YC(w_mem_inst_add_2_root_add_945_3_carry[29]), .YS(w_mem_inst_N668));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_29 ( .A(w_mem_inst_N610),  .B(w_mem_inst_w_mem[221]),  .C(w_mem_inst_add_2_root_add_945_3_carry[29]), .YC(w_mem_inst_add_2_root_add_945_3_carry[30]), .YS(w_mem_inst_N669));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_30 ( .A(w_mem_inst_N609),  .B(w_mem_inst_w_mem[222]),  .C(w_mem_inst_add_2_root_add_945_3_carry[30]), .YC(w_mem_inst_add_2_root_add_945_3_carry[31]), .YS(w_mem_inst_N670));
   FAX1 w_mem_inst_add_2_root_add_945_3_U1_31 ( .A(w_mem_inst_N608),  .B(w_mem_inst_w_mem[223]),  .C(w_mem_inst_add_2_root_add_945_3_carry[31]), .YS(w_mem_inst_N671));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_1 ( .A(w_mem_inst_N606),  .B(w_mem_inst_w_mem[481]),  .C(n2965), .YC(w_mem_inst_add_1_root_add_945_3_carry[2]), .YS(w_mem_inst_N673));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_2 ( .A(w_mem_inst_N605),  .B(w_mem_inst_w_mem[482]),  .C(w_mem_inst_add_1_root_add_945_3_carry[2]), .YC(w_mem_inst_add_1_root_add_945_3_carry[3]), .YS(w_mem_inst_N674));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_3 ( .A(w_mem_inst_N604),  .B(w_mem_inst_w_mem[483]),  .C(w_mem_inst_add_1_root_add_945_3_carry[3]), .YC(w_mem_inst_add_1_root_add_945_3_carry[4]), .YS(w_mem_inst_N675));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_4 ( .A(w_mem_inst_N603),  .B(w_mem_inst_w_mem[484]),  .C(w_mem_inst_add_1_root_add_945_3_carry[4]), .YC(w_mem_inst_add_1_root_add_945_3_carry[5]), .YS(w_mem_inst_N676));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_5 ( .A(w_mem_inst_N602),  .B(w_mem_inst_w_mem[485]),  .C(w_mem_inst_add_1_root_add_945_3_carry[5]), .YC(w_mem_inst_add_1_root_add_945_3_carry[6]), .YS(w_mem_inst_N677));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_6 ( .A(w_mem_inst_N601),  .B(w_mem_inst_w_mem[486]),  .C(w_mem_inst_add_1_root_add_945_3_carry[6]), .YC(w_mem_inst_add_1_root_add_945_3_carry[7]), .YS(w_mem_inst_N678));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_7 ( .A(w_mem_inst_N600),  .B(w_mem_inst_w_mem[487]),  .C(w_mem_inst_add_1_root_add_945_3_carry[7]), .YC(w_mem_inst_add_1_root_add_945_3_carry[8]), .YS(w_mem_inst_N679));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_8 ( .A(w_mem_inst_N599),  .B(w_mem_inst_w_mem[488]),  .C(w_mem_inst_add_1_root_add_945_3_carry[8]), .YC(w_mem_inst_add_1_root_add_945_3_carry[9]), .YS(w_mem_inst_N680));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_9 ( .A(w_mem_inst_N598),  .B(w_mem_inst_w_mem[489]),  .C(w_mem_inst_add_1_root_add_945_3_carry[9]), .YC(w_mem_inst_add_1_root_add_945_3_carry[10]), .YS(w_mem_inst_N681));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_10 ( .A(w_mem_inst_N597),  .B(w_mem_inst_w_mem[490]),  .C(w_mem_inst_add_1_root_add_945_3_carry[10]), .YC(w_mem_inst_add_1_root_add_945_3_carry[11]), .YS(w_mem_inst_N682));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_11 ( .A(w_mem_inst_N596),  .B(w_mem_inst_w_mem[491]),  .C(w_mem_inst_add_1_root_add_945_3_carry[11]), .YC(w_mem_inst_add_1_root_add_945_3_carry[12]), .YS(w_mem_inst_N683));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_12 ( .A(w_mem_inst_N595),  .B(w_mem_inst_w_mem[492]),  .C(w_mem_inst_add_1_root_add_945_3_carry[12]), .YC(w_mem_inst_add_1_root_add_945_3_carry[13]), .YS(w_mem_inst_N684));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_13 ( .A(w_mem_inst_N594),  .B(w_mem_inst_w_mem[493]),  .C(w_mem_inst_add_1_root_add_945_3_carry[13]), .YC(w_mem_inst_add_1_root_add_945_3_carry[14]), .YS(w_mem_inst_N685));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_14 ( .A(w_mem_inst_N593),  .B(w_mem_inst_w_mem[494]),  .C(w_mem_inst_add_1_root_add_945_3_carry[14]), .YC(w_mem_inst_add_1_root_add_945_3_carry[15]), .YS(w_mem_inst_N686));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_15 ( .A(w_mem_inst_N592),  .B(w_mem_inst_w_mem[495]),  .C(w_mem_inst_add_1_root_add_945_3_carry[15]), .YC(w_mem_inst_add_1_root_add_945_3_carry[16]), .YS(w_mem_inst_N687));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_16 ( .A(w_mem_inst_N591),  .B(w_mem_inst_w_mem[496]),  .C(w_mem_inst_add_1_root_add_945_3_carry[16]), .YC(w_mem_inst_add_1_root_add_945_3_carry[17]), .YS(w_mem_inst_N688));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_17 ( .A(w_mem_inst_N590),  .B(w_mem_inst_w_mem[497]),  .C(w_mem_inst_add_1_root_add_945_3_carry[17]), .YC(w_mem_inst_add_1_root_add_945_3_carry[18]), .YS(w_mem_inst_N689));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_18 ( .A(w_mem_inst_N589),  .B(w_mem_inst_w_mem[498]),  .C(w_mem_inst_add_1_root_add_945_3_carry[18]), .YC(w_mem_inst_add_1_root_add_945_3_carry[19]), .YS(w_mem_inst_N690));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_19 ( .A(w_mem_inst_N588),  .B(w_mem_inst_w_mem[499]),  .C(w_mem_inst_add_1_root_add_945_3_carry[19]), .YC(w_mem_inst_add_1_root_add_945_3_carry[20]), .YS(w_mem_inst_N691));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_20 ( .A(w_mem_inst_N587),  .B(w_mem_inst_w_mem[500]),  .C(w_mem_inst_add_1_root_add_945_3_carry[20]), .YC(w_mem_inst_add_1_root_add_945_3_carry[21]), .YS(w_mem_inst_N692));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_21 ( .A(w_mem_inst_N586),  .B(w_mem_inst_w_mem[501]),  .C(w_mem_inst_add_1_root_add_945_3_carry[21]), .YC(w_mem_inst_add_1_root_add_945_3_carry[22]), .YS(w_mem_inst_N693));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_22 ( .A(w_mem_inst_N585),  .B(w_mem_inst_w_mem[502]),  .C(w_mem_inst_add_1_root_add_945_3_carry[22]), .YC(w_mem_inst_add_1_root_add_945_3_carry[23]), .YS(w_mem_inst_N694));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_23 ( .A(w_mem_inst_N584),  .B(w_mem_inst_w_mem[503]),  .C(w_mem_inst_add_1_root_add_945_3_carry[23]), .YC(w_mem_inst_add_1_root_add_945_3_carry[24]), .YS(w_mem_inst_N695));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_24 ( .A(w_mem_inst_N583),  .B(w_mem_inst_w_mem[504]),  .C(w_mem_inst_add_1_root_add_945_3_carry[24]), .YC(w_mem_inst_add_1_root_add_945_3_carry[25]), .YS(w_mem_inst_N696));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_25 ( .A(w_mem_inst_N582),  .B(w_mem_inst_w_mem[505]),  .C(w_mem_inst_add_1_root_add_945_3_carry[25]), .YC(w_mem_inst_add_1_root_add_945_3_carry[26]), .YS(w_mem_inst_N697));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_26 ( .A(w_mem_inst_N581),  .B(w_mem_inst_w_mem[506]),  .C(w_mem_inst_add_1_root_add_945_3_carry[26]), .YC(w_mem_inst_add_1_root_add_945_3_carry[27]), .YS(w_mem_inst_N698));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_27 ( .A(w_mem_inst_N580),  .B(w_mem_inst_w_mem[507]),  .C(w_mem_inst_add_1_root_add_945_3_carry[27]), .YC(w_mem_inst_add_1_root_add_945_3_carry[28]), .YS(w_mem_inst_N699));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_28 ( .A(w_mem_inst_N579),  .B(w_mem_inst_w_mem[508]),  .C(w_mem_inst_add_1_root_add_945_3_carry[28]), .YC(w_mem_inst_add_1_root_add_945_3_carry[29]), .YS(w_mem_inst_N700));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_29 ( .A(w_mem_inst_N578),  .B(w_mem_inst_w_mem[509]),  .C(w_mem_inst_add_1_root_add_945_3_carry[29]), .YC(w_mem_inst_add_1_root_add_945_3_carry[30]), .YS(w_mem_inst_N701));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_30 ( .A(w_mem_inst_N577),  .B(w_mem_inst_w_mem[510]),  .C(w_mem_inst_add_1_root_add_945_3_carry[30]), .YC(w_mem_inst_add_1_root_add_945_3_carry[31]), .YS(w_mem_inst_N702));
   FAX1 w_mem_inst_add_1_root_add_945_3_U1_31 ( .A(w_mem_inst_N576),  .B(w_mem_inst_w_mem[511]),  .C(w_mem_inst_add_1_root_add_945_3_carry[31]), .YS(w_mem_inst_N703));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_1 ( .A(w_mem_inst_N641),  .B(w_mem_inst_N673),  .C(n2962), .YC(w_mem_inst_add_0_root_add_945_3_carry[2]), .YS(w_mem_inst_w_new[1]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_2 ( .A(w_mem_inst_N642),  .B(w_mem_inst_N674),  .C(w_mem_inst_add_0_root_add_945_3_carry[2]), .YC(w_mem_inst_add_0_root_add_945_3_carry[3]), .YS(w_mem_inst_w_new[2]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_3 ( .A(w_mem_inst_N643),  .B(w_mem_inst_N675),  .C(w_mem_inst_add_0_root_add_945_3_carry[3]), .YC(w_mem_inst_add_0_root_add_945_3_carry[4]), .YS(w_mem_inst_w_new[3]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_4 ( .A(w_mem_inst_N644),  .B(w_mem_inst_N676),  .C(w_mem_inst_add_0_root_add_945_3_carry[4]), .YC(w_mem_inst_add_0_root_add_945_3_carry[5]), .YS(w_mem_inst_w_new[4]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_5 ( .A(w_mem_inst_N645),  .B(w_mem_inst_N677),  .C(w_mem_inst_add_0_root_add_945_3_carry[5]), .YC(w_mem_inst_add_0_root_add_945_3_carry[6]), .YS(w_mem_inst_w_new[5]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_6 ( .A(w_mem_inst_N646),  .B(w_mem_inst_N678),  .C(w_mem_inst_add_0_root_add_945_3_carry[6]), .YC(w_mem_inst_add_0_root_add_945_3_carry[7]), .YS(w_mem_inst_w_new[6]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_7 ( .A(w_mem_inst_N647),  .B(w_mem_inst_N679),  .C(w_mem_inst_add_0_root_add_945_3_carry[7]), .YC(w_mem_inst_add_0_root_add_945_3_carry[8]), .YS(w_mem_inst_w_new[7]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_8 ( .A(w_mem_inst_N648),  .B(w_mem_inst_N680),  .C(w_mem_inst_add_0_root_add_945_3_carry[8]), .YC(w_mem_inst_add_0_root_add_945_3_carry[9]), .YS(w_mem_inst_w_new[8]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_9 ( .A(w_mem_inst_N649),  .B(w_mem_inst_N681),  .C(w_mem_inst_add_0_root_add_945_3_carry[9]), .YC(w_mem_inst_add_0_root_add_945_3_carry[10]), .YS(w_mem_inst_w_new[9]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_10 ( .A(w_mem_inst_N650),  .B(w_mem_inst_N682),  .C(w_mem_inst_add_0_root_add_945_3_carry[10]), .YC(w_mem_inst_add_0_root_add_945_3_carry[11]), .YS(w_mem_inst_w_new[10]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_11 ( .A(w_mem_inst_N651),  .B(w_mem_inst_N683),  .C(w_mem_inst_add_0_root_add_945_3_carry[11]), .YC(w_mem_inst_add_0_root_add_945_3_carry[12]), .YS(w_mem_inst_w_new[11]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_12 ( .A(w_mem_inst_N652),  .B(w_mem_inst_N684),  .C(w_mem_inst_add_0_root_add_945_3_carry[12]), .YC(w_mem_inst_add_0_root_add_945_3_carry[13]), .YS(w_mem_inst_w_new[12]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_13 ( .A(w_mem_inst_N653),  .B(w_mem_inst_N685),  .C(w_mem_inst_add_0_root_add_945_3_carry[13]), .YC(w_mem_inst_add_0_root_add_945_3_carry[14]), .YS(w_mem_inst_w_new[13]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_14 ( .A(w_mem_inst_N654),  .B(w_mem_inst_N686),  .C(w_mem_inst_add_0_root_add_945_3_carry[14]), .YC(w_mem_inst_add_0_root_add_945_3_carry[15]), .YS(w_mem_inst_w_new[14]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_15 ( .A(w_mem_inst_N655),  .B(w_mem_inst_N687),  .C(w_mem_inst_add_0_root_add_945_3_carry[15]), .YC(w_mem_inst_add_0_root_add_945_3_carry[16]), .YS(w_mem_inst_w_new[15]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_16 ( .A(w_mem_inst_N656),  .B(w_mem_inst_N688),  .C(w_mem_inst_add_0_root_add_945_3_carry[16]), .YC(w_mem_inst_add_0_root_add_945_3_carry[17]), .YS(w_mem_inst_w_new[16]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_17 ( .A(w_mem_inst_N657),  .B(w_mem_inst_N689),  .C(w_mem_inst_add_0_root_add_945_3_carry[17]), .YC(w_mem_inst_add_0_root_add_945_3_carry[18]), .YS(w_mem_inst_w_new[17]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_18 ( .A(w_mem_inst_N658),  .B(w_mem_inst_N690),  .C(w_mem_inst_add_0_root_add_945_3_carry[18]), .YC(w_mem_inst_add_0_root_add_945_3_carry[19]), .YS(w_mem_inst_w_new[18]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_19 ( .A(w_mem_inst_N659),  .B(w_mem_inst_N691),  .C(w_mem_inst_add_0_root_add_945_3_carry[19]), .YC(w_mem_inst_add_0_root_add_945_3_carry[20]), .YS(w_mem_inst_w_new[19]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_20 ( .A(w_mem_inst_N660),  .B(w_mem_inst_N692),  .C(w_mem_inst_add_0_root_add_945_3_carry[20]), .YC(w_mem_inst_add_0_root_add_945_3_carry[21]), .YS(w_mem_inst_w_new[20]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_21 ( .A(w_mem_inst_N661),  .B(w_mem_inst_N693),  .C(w_mem_inst_add_0_root_add_945_3_carry[21]), .YC(w_mem_inst_add_0_root_add_945_3_carry[22]), .YS(w_mem_inst_w_new[21]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_22 ( .A(w_mem_inst_N662),  .B(w_mem_inst_N694),  .C(w_mem_inst_add_0_root_add_945_3_carry[22]), .YC(w_mem_inst_add_0_root_add_945_3_carry[23]), .YS(w_mem_inst_w_new[22]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_23 ( .A(w_mem_inst_N663),  .B(w_mem_inst_N695),  .C(w_mem_inst_add_0_root_add_945_3_carry[23]), .YC(w_mem_inst_add_0_root_add_945_3_carry[24]), .YS(w_mem_inst_w_new[23]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_24 ( .A(w_mem_inst_N664),  .B(w_mem_inst_N696),  .C(w_mem_inst_add_0_root_add_945_3_carry[24]), .YC(w_mem_inst_add_0_root_add_945_3_carry[25]), .YS(w_mem_inst_w_new[24]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_25 ( .A(w_mem_inst_N665),  .B(w_mem_inst_N697),  .C(w_mem_inst_add_0_root_add_945_3_carry[25]), .YC(w_mem_inst_add_0_root_add_945_3_carry[26]), .YS(w_mem_inst_w_new[25]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_26 ( .A(w_mem_inst_N666),  .B(w_mem_inst_N698),  .C(w_mem_inst_add_0_root_add_945_3_carry[26]), .YC(w_mem_inst_add_0_root_add_945_3_carry[27]), .YS(w_mem_inst_w_new[26]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_27 ( .A(w_mem_inst_N667),  .B(w_mem_inst_N699),  .C(w_mem_inst_add_0_root_add_945_3_carry[27]), .YC(w_mem_inst_add_0_root_add_945_3_carry[28]), .YS(w_mem_inst_w_new[27]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_28 ( .A(w_mem_inst_N668),  .B(w_mem_inst_N700),  .C(w_mem_inst_add_0_root_add_945_3_carry[28]), .YC(w_mem_inst_add_0_root_add_945_3_carry[29]), .YS(w_mem_inst_w_new[28]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_29 ( .A(w_mem_inst_N669),  .B(w_mem_inst_N701),  .C(w_mem_inst_add_0_root_add_945_3_carry[29]), .YC(w_mem_inst_add_0_root_add_945_3_carry[30]), .YS(w_mem_inst_w_new[29]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_30 ( .A(w_mem_inst_N670),  .B(w_mem_inst_N702),  .C(w_mem_inst_add_0_root_add_945_3_carry[30]), .YC(w_mem_inst_add_0_root_add_945_3_carry[31]), .YS(w_mem_inst_w_new[30]));
   FAX1 w_mem_inst_add_0_root_add_945_3_U1_31 ( .A(w_mem_inst_N671),  .B(w_mem_inst_N703),  .C(w_mem_inst_add_0_root_add_945_3_carry[31]), .YS(w_mem_inst_w_new[31]));
   HAX1 w_mem_inst_add_1008_U1_1_1 ( .A(w_mem_inst_w_ctr_reg[1]),  .B(w_mem_inst_w_ctr_reg[0]), .YC(w_mem_inst_add_1008_carry[2]), .YS(w_mem_inst_N711));
   HAX1 w_mem_inst_add_1008_U1_1_2 ( .A(w_mem_inst_w_ctr_reg[2]),  .B(w_mem_inst_add_1008_carry[2]), .YC(w_mem_inst_add_1008_carry[3]), .YS(w_mem_inst_N712));
   HAX1 w_mem_inst_add_1008_U1_1_3 ( .A(w_mem_inst_w_ctr_reg[3]),  .B(w_mem_inst_add_1008_carry[3]), .YC(w_mem_inst_add_1008_carry[4]), .YS(w_mem_inst_N713));
   HAX1 w_mem_inst_add_1008_U1_1_4 ( .A(w_mem_inst_w_ctr_reg[4]),  .B(w_mem_inst_add_1008_carry[4]), .YC(w_mem_inst_add_1008_carry[5]), .YS(w_mem_inst_N714));
   HAX1 add_420_U1_1_1 ( .A(t_ctr_reg[1]),  .B(t_ctr_reg[0]), .YC(add_420_carry[2]), .YS(N1615));
   HAX1 add_420_U1_1_2 ( .A(t_ctr_reg[2]),  .B(add_420_carry[2]), .YC(add_420_carry[3]), .YS(N1616));
   HAX1 add_420_U1_1_3 ( .A(t_ctr_reg[3]),  .B(add_420_carry[3]), .YC(add_420_carry[4]), .YS(N1617));
   HAX1 add_420_U1_1_4 ( .A(t_ctr_reg[4]),  .B(add_420_carry[4]), .YC(add_420_carry[5]), .YS(N1618));
   FAX1 add_392_U1_1 ( .A(d_reg[1]),  .B(t1[1]),  .C(n2967), .YC(add_392_carry[2]), .YS(N1580));
   FAX1 add_392_U1_2 ( .A(d_reg[2]),  .B(t1[2]),  .C(add_392_carry[2]), .YC(add_392_carry[3]), .YS(N1581));
   FAX1 add_392_U1_3 ( .A(d_reg[3]),  .B(t1[3]),  .C(add_392_carry[3]), .YC(add_392_carry[4]), .YS(N1582));
   FAX1 add_392_U1_4 ( .A(d_reg[4]),  .B(t1[4]),  .C(add_392_carry[4]), .YC(add_392_carry[5]), .YS(N1583));
   FAX1 add_392_U1_5 ( .A(d_reg[5]),  .B(t1[5]),  .C(add_392_carry[5]), .YC(add_392_carry[6]), .YS(N1584));
   FAX1 add_392_U1_6 ( .A(d_reg[6]),  .B(t1[6]),  .C(add_392_carry[6]), .YC(add_392_carry[7]), .YS(N1585));
   FAX1 add_392_U1_7 ( .A(d_reg[7]),  .B(t1[7]),  .C(add_392_carry[7]), .YC(add_392_carry[8]), .YS(N1586));
   FAX1 add_392_U1_8 ( .A(d_reg[8]),  .B(t1[8]),  .C(add_392_carry[8]), .YC(add_392_carry[9]), .YS(N1587));
   FAX1 add_392_U1_9 ( .A(d_reg[9]),  .B(t1[9]),  .C(add_392_carry[9]), .YC(add_392_carry[10]), .YS(N1588));
   FAX1 add_392_U1_10 ( .A(d_reg[10]),  .B(t1[10]),  .C(add_392_carry[10]), .YC(add_392_carry[11]), .YS(N1589));
   FAX1 add_392_U1_11 ( .A(d_reg[11]),  .B(t1[11]),  .C(add_392_carry[11]), .YC(add_392_carry[12]), .YS(N1590));
   FAX1 add_392_U1_12 ( .A(d_reg[12]),  .B(t1[12]),  .C(add_392_carry[12]), .YC(add_392_carry[13]), .YS(N1591));
   FAX1 add_392_U1_13 ( .A(d_reg[13]),  .B(t1[13]),  .C(add_392_carry[13]), .YC(add_392_carry[14]), .YS(N1592));
   FAX1 add_392_U1_14 ( .A(d_reg[14]),  .B(t1[14]),  .C(add_392_carry[14]), .YC(add_392_carry[15]), .YS(N1593));
   FAX1 add_392_U1_15 ( .A(d_reg[15]),  .B(t1[15]),  .C(add_392_carry[15]), .YC(add_392_carry[16]), .YS(N1594));
   FAX1 add_392_U1_16 ( .A(d_reg[16]),  .B(t1[16]),  .C(add_392_carry[16]), .YC(add_392_carry[17]), .YS(N1595));
   FAX1 add_392_U1_17 ( .A(d_reg[17]),  .B(t1[17]),  .C(add_392_carry[17]), .YC(add_392_carry[18]), .YS(N1596));
   FAX1 add_392_U1_18 ( .A(d_reg[18]),  .B(t1[18]),  .C(add_392_carry[18]), .YC(add_392_carry[19]), .YS(N1597));
   FAX1 add_392_U1_19 ( .A(d_reg[19]),  .B(t1[19]),  .C(add_392_carry[19]), .YC(add_392_carry[20]), .YS(N1598));
   FAX1 add_392_U1_20 ( .A(d_reg[20]),  .B(t1[20]),  .C(add_392_carry[20]), .YC(add_392_carry[21]), .YS(N1599));
   FAX1 add_392_U1_21 ( .A(d_reg[21]),  .B(t1[21]),  .C(add_392_carry[21]), .YC(add_392_carry[22]), .YS(N1600));
   FAX1 add_392_U1_22 ( .A(d_reg[22]),  .B(t1[22]),  .C(add_392_carry[22]), .YC(add_392_carry[23]), .YS(N1601));
   FAX1 add_392_U1_23 ( .A(d_reg[23]),  .B(t1[23]),  .C(add_392_carry[23]), .YC(add_392_carry[24]), .YS(N1602));
   FAX1 add_392_U1_24 ( .A(d_reg[24]),  .B(t1[24]),  .C(add_392_carry[24]), .YC(add_392_carry[25]), .YS(N1603));
   FAX1 add_392_U1_25 ( .A(d_reg[25]),  .B(t1[25]),  .C(add_392_carry[25]), .YC(add_392_carry[26]), .YS(N1604));
   FAX1 add_392_U1_26 ( .A(d_reg[26]),  .B(t1[26]),  .C(add_392_carry[26]), .YC(add_392_carry[27]), .YS(N1605));
   FAX1 add_392_U1_27 ( .A(d_reg[27]),  .B(t1[27]),  .C(add_392_carry[27]), .YC(add_392_carry[28]), .YS(N1606));
   FAX1 add_392_U1_28 ( .A(d_reg[28]),  .B(t1[28]),  .C(add_392_carry[28]), .YC(add_392_carry[29]), .YS(N1607));
   FAX1 add_392_U1_29 ( .A(d_reg[29]),  .B(t1[29]),  .C(add_392_carry[29]), .YC(add_392_carry[30]), .YS(N1608));
   FAX1 add_392_U1_30 ( .A(d_reg[30]),  .B(t1[30]),  .C(add_392_carry[30]), .YC(add_392_carry[31]), .YS(N1609));
   FAX1 add_392_U1_31 ( .A(d_reg[31]),  .B(t1[31]),  .C(add_392_carry[31]), .YS(N1610));
   FAX1 add_0_root_add_388_U1_1 ( .A(N1028),  .B(t2[1]),  .C(n2960), .YC(add_0_root_add_388_carry[2]), .YS(N1548));
   FAX1 add_0_root_add_388_U1_2 ( .A(n6194),  .B(t2[2]),  .C(add_0_root_add_388_carry[2]), .YC(add_0_root_add_388_carry[3]), .YS(N1549));
   FAX1 add_0_root_add_388_U1_3 ( .A(N1026),  .B(t2[3]),  .C(add_0_root_add_388_carry[3]), .YC(add_0_root_add_388_carry[4]), .YS(N1550));
   FAX1 add_0_root_add_388_U1_4 ( .A(N1025),  .B(t2[4]),  .C(add_0_root_add_388_carry[4]), .YC(add_0_root_add_388_carry[5]), .YS(N1551));
   FAX1 add_0_root_add_388_U1_5 ( .A(N1024),  .B(t2[5]),  .C(add_0_root_add_388_carry[5]), .YC(add_0_root_add_388_carry[6]), .YS(N1552));
   FAX1 add_0_root_add_388_U1_6 ( .A(N1023),  .B(t2[6]),  .C(add_0_root_add_388_carry[6]), .YC(add_0_root_add_388_carry[7]), .YS(N1553));
   FAX1 add_0_root_add_388_U1_7 ( .A(N1022),  .B(t2[7]),  .C(add_0_root_add_388_carry[7]), .YC(add_0_root_add_388_carry[8]), .YS(N1554));
   FAX1 add_0_root_add_388_U1_8 ( .A(N1021),  .B(t2[8]),  .C(add_0_root_add_388_carry[8]), .YC(add_0_root_add_388_carry[9]), .YS(N1555));
   FAX1 add_0_root_add_388_U1_9 ( .A(n6195),  .B(t2[9]),  .C(add_0_root_add_388_carry[9]), .YC(add_0_root_add_388_carry[10]), .YS(N1556));
   FAX1 add_0_root_add_388_U1_10 ( .A(n6196),  .B(t2[10]),  .C(add_0_root_add_388_carry[10]), .YC(add_0_root_add_388_carry[11]), .YS(N1557));
   FAX1 add_0_root_add_388_U1_11 ( .A(N1018),  .B(t2[11]),  .C(add_0_root_add_388_carry[11]), .YC(add_0_root_add_388_carry[12]), .YS(N1558));
   FAX1 add_0_root_add_388_U1_12 ( .A(N1017),  .B(t2[12]),  .C(add_0_root_add_388_carry[12]), .YC(add_0_root_add_388_carry[13]), .YS(N1559));
   FAX1 add_0_root_add_388_U1_13 ( .A(N1016),  .B(t2[13]),  .C(add_0_root_add_388_carry[13]), .YC(add_0_root_add_388_carry[14]), .YS(N1560));
   FAX1 add_0_root_add_388_U1_14 ( .A(N1015),  .B(t2[14]),  .C(add_0_root_add_388_carry[14]), .YC(add_0_root_add_388_carry[15]), .YS(N1561));
   FAX1 add_0_root_add_388_U1_15 ( .A(N1014),  .B(t2[15]),  .C(add_0_root_add_388_carry[15]), .YC(add_0_root_add_388_carry[16]), .YS(N1562));
   FAX1 add_0_root_add_388_U1_16 ( .A(N1013),  .B(t2[16]),  .C(add_0_root_add_388_carry[16]), .YC(add_0_root_add_388_carry[17]), .YS(N1563));
   FAX1 add_0_root_add_388_U1_17 ( .A(N1012),  .B(t2[17]),  .C(add_0_root_add_388_carry[17]), .YC(add_0_root_add_388_carry[18]), .YS(N1564));
   FAX1 add_0_root_add_388_U1_18 ( .A(N1011),  .B(t2[18]),  .C(add_0_root_add_388_carry[18]), .YC(add_0_root_add_388_carry[19]), .YS(N1565));
   FAX1 add_0_root_add_388_U1_19 ( .A(N1010),  .B(t2[19]),  .C(add_0_root_add_388_carry[19]), .YC(add_0_root_add_388_carry[20]), .YS(N1566));
   FAX1 add_0_root_add_388_U1_20 ( .A(N1009),  .B(t2[20]),  .C(add_0_root_add_388_carry[20]), .YC(add_0_root_add_388_carry[21]), .YS(N1567));
   FAX1 add_0_root_add_388_U1_21 ( .A(N1008),  .B(t2[21]),  .C(add_0_root_add_388_carry[21]), .YC(add_0_root_add_388_carry[22]), .YS(N1568));
   FAX1 add_0_root_add_388_U1_22 ( .A(N1007),  .B(t2[22]),  .C(add_0_root_add_388_carry[22]), .YC(add_0_root_add_388_carry[23]), .YS(N1569));
   FAX1 add_0_root_add_388_U1_23 ( .A(N1006),  .B(t2[23]),  .C(add_0_root_add_388_carry[23]), .YC(add_0_root_add_388_carry[24]), .YS(N1570));
   FAX1 add_0_root_add_388_U1_24 ( .A(N1005),  .B(t2[24]),  .C(add_0_root_add_388_carry[24]), .YC(add_0_root_add_388_carry[25]), .YS(N1571));
   FAX1 add_0_root_add_388_U1_25 ( .A(n6197),  .B(t2[25]),  .C(add_0_root_add_388_carry[25]), .YC(add_0_root_add_388_carry[26]), .YS(N1572));
   FAX1 add_0_root_add_388_U1_26 ( .A(N1003),  .B(t2[26]),  .C(add_0_root_add_388_carry[26]), .YC(add_0_root_add_388_carry[27]), .YS(N1573));
   FAX1 add_0_root_add_388_U1_27 ( .A(n6198),  .B(t2[27]),  .C(add_0_root_add_388_carry[27]), .YC(add_0_root_add_388_carry[28]), .YS(N1574));
   FAX1 add_0_root_add_388_U1_28 ( .A(N1001),  .B(t2[28]),  .C(add_0_root_add_388_carry[28]), .YC(add_0_root_add_388_carry[29]), .YS(N1575));
   FAX1 add_0_root_add_388_U1_29 ( .A(n6199),  .B(t2[29]),  .C(add_0_root_add_388_carry[29]), .YC(add_0_root_add_388_carry[30]), .YS(N1576));
   FAX1 add_0_root_add_388_U1_30 ( .A(N999),  .B(t2[30]),  .C(add_0_root_add_388_carry[30]), .YC(add_0_root_add_388_carry[31]), .YS(N1577));
   FAX1 add_0_root_add_388_U1_31 ( .A(N998),  .B(t2[31]),  .C(add_0_root_add_388_carry[31]), .YS(N1578));
   FAX1 add_1_root_add_388_U1_1 ( .A(t1[1]),  .B(N996),  .C(n2963), .YC(add_1_root_add_388_carry[2]), .YS(t2[1]));
   FAX1 add_1_root_add_388_U1_2 ( .A(t1[2]),  .B(N995),  .C(add_1_root_add_388_carry[2]), .YC(add_1_root_add_388_carry[3]), .YS(t2[2]));
   FAX1 add_1_root_add_388_U1_3 ( .A(t1[3]),  .B(N994),  .C(add_1_root_add_388_carry[3]), .YC(add_1_root_add_388_carry[4]), .YS(t2[3]));
   FAX1 add_1_root_add_388_U1_4 ( .A(t1[4]),  .B(N993),  .C(add_1_root_add_388_carry[4]), .YC(add_1_root_add_388_carry[5]), .YS(t2[4]));
   FAX1 add_1_root_add_388_U1_5 ( .A(t1[5]),  .B(N992),  .C(add_1_root_add_388_carry[5]), .YC(add_1_root_add_388_carry[6]), .YS(t2[5]));
   FAX1 add_1_root_add_388_U1_6 ( .A(t1[6]),  .B(N991),  .C(add_1_root_add_388_carry[6]), .YC(add_1_root_add_388_carry[7]), .YS(t2[6]));
   FAX1 add_1_root_add_388_U1_7 ( .A(t1[7]),  .B(N990),  .C(add_1_root_add_388_carry[7]), .YC(add_1_root_add_388_carry[8]), .YS(t2[7]));
   FAX1 add_1_root_add_388_U1_8 ( .A(t1[8]),  .B(N989),  .C(add_1_root_add_388_carry[8]), .YC(add_1_root_add_388_carry[9]), .YS(t2[8]));
   FAX1 add_1_root_add_388_U1_9 ( .A(t1[9]),  .B(N988),  .C(add_1_root_add_388_carry[9]), .YC(add_1_root_add_388_carry[10]), .YS(t2[9]));
   FAX1 add_1_root_add_388_U1_10 ( .A(t1[10]),  .B(N987),  .C(add_1_root_add_388_carry[10]), .YC(add_1_root_add_388_carry[11]), .YS(t2[10]));
   FAX1 add_1_root_add_388_U1_11 ( .A(t1[11]),  .B(N986),  .C(add_1_root_add_388_carry[11]), .YC(add_1_root_add_388_carry[12]), .YS(t2[11]));
   FAX1 add_1_root_add_388_U1_12 ( .A(t1[12]),  .B(N985),  .C(add_1_root_add_388_carry[12]), .YC(add_1_root_add_388_carry[13]), .YS(t2[12]));
   FAX1 add_1_root_add_388_U1_13 ( .A(t1[13]),  .B(N984),  .C(add_1_root_add_388_carry[13]), .YC(add_1_root_add_388_carry[14]), .YS(t2[13]));
   FAX1 add_1_root_add_388_U1_14 ( .A(t1[14]),  .B(N983),  .C(add_1_root_add_388_carry[14]), .YC(add_1_root_add_388_carry[15]), .YS(t2[14]));
   FAX1 add_1_root_add_388_U1_15 ( .A(t1[15]),  .B(N982),  .C(add_1_root_add_388_carry[15]), .YC(add_1_root_add_388_carry[16]), .YS(t2[15]));
   FAX1 add_1_root_add_388_U1_16 ( .A(t1[16]),  .B(N981),  .C(add_1_root_add_388_carry[16]), .YC(add_1_root_add_388_carry[17]), .YS(t2[16]));
   FAX1 add_1_root_add_388_U1_17 ( .A(t1[17]),  .B(N980),  .C(add_1_root_add_388_carry[17]), .YC(add_1_root_add_388_carry[18]), .YS(t2[17]));
   FAX1 add_1_root_add_388_U1_18 ( .A(t1[18]),  .B(N979),  .C(add_1_root_add_388_carry[18]), .YC(add_1_root_add_388_carry[19]), .YS(t2[18]));
   FAX1 add_1_root_add_388_U1_19 ( .A(t1[19]),  .B(N978),  .C(add_1_root_add_388_carry[19]), .YC(add_1_root_add_388_carry[20]), .YS(t2[19]));
   FAX1 add_1_root_add_388_U1_20 ( .A(t1[20]),  .B(N977),  .C(add_1_root_add_388_carry[20]), .YC(add_1_root_add_388_carry[21]), .YS(t2[20]));
   FAX1 add_1_root_add_388_U1_21 ( .A(t1[21]),  .B(N976),  .C(add_1_root_add_388_carry[21]), .YC(add_1_root_add_388_carry[22]), .YS(t2[21]));
   FAX1 add_1_root_add_388_U1_22 ( .A(t1[22]),  .B(N975),  .C(add_1_root_add_388_carry[22]), .YC(add_1_root_add_388_carry[23]), .YS(t2[22]));
   FAX1 add_1_root_add_388_U1_23 ( .A(t1[23]),  .B(N974),  .C(add_1_root_add_388_carry[23]), .YC(add_1_root_add_388_carry[24]), .YS(t2[23]));
   FAX1 add_1_root_add_388_U1_24 ( .A(t1[24]),  .B(N973),  .C(add_1_root_add_388_carry[24]), .YC(add_1_root_add_388_carry[25]), .YS(t2[24]));
   FAX1 add_1_root_add_388_U1_25 ( .A(t1[25]),  .B(N972),  .C(add_1_root_add_388_carry[25]), .YC(add_1_root_add_388_carry[26]), .YS(t2[25]));
   FAX1 add_1_root_add_388_U1_26 ( .A(t1[26]),  .B(N971),  .C(add_1_root_add_388_carry[26]), .YC(add_1_root_add_388_carry[27]), .YS(t2[26]));
   FAX1 add_1_root_add_388_U1_27 ( .A(t1[27]),  .B(N970),  .C(add_1_root_add_388_carry[27]), .YC(add_1_root_add_388_carry[28]), .YS(t2[27]));
   FAX1 add_1_root_add_388_U1_28 ( .A(t1[28]),  .B(N969),  .C(add_1_root_add_388_carry[28]), .YC(add_1_root_add_388_carry[29]), .YS(t2[28]));
   FAX1 add_1_root_add_388_U1_29 ( .A(t1[29]),  .B(N968),  .C(add_1_root_add_388_carry[29]), .YC(add_1_root_add_388_carry[30]), .YS(t2[29]));
   FAX1 add_1_root_add_388_U1_30 ( .A(t1[30]),  .B(N967),  .C(add_1_root_add_388_carry[30]), .YC(add_1_root_add_388_carry[31]), .YS(t2[30]));
   FAX1 add_1_root_add_388_U1_31 ( .A(t1[31]),  .B(N966),  .C(add_1_root_add_388_carry[31]), .YS(t2[31]));
   FAX1 add_0_root_add_317_4_U1_1 ( .A(N903),  .B(N935),  .C(n2959), .YC(add_0_root_add_317_4_carry[2]), .YS(t1[1]));
   FAX1 add_0_root_add_317_4_U1_2 ( .A(N904),  .B(N936),  .C(add_0_root_add_317_4_carry[2]), .YC(add_0_root_add_317_4_carry[3]), .YS(t1[2]));
   FAX1 add_0_root_add_317_4_U1_3 ( .A(N905),  .B(N937),  .C(add_0_root_add_317_4_carry[3]), .YC(add_0_root_add_317_4_carry[4]), .YS(t1[3]));
   FAX1 add_0_root_add_317_4_U1_4 ( .A(N906),  .B(N938),  .C(add_0_root_add_317_4_carry[4]), .YC(add_0_root_add_317_4_carry[5]), .YS(t1[4]));
   FAX1 add_0_root_add_317_4_U1_5 ( .A(N907),  .B(N939),  .C(add_0_root_add_317_4_carry[5]), .YC(add_0_root_add_317_4_carry[6]), .YS(t1[5]));
   FAX1 add_0_root_add_317_4_U1_6 ( .A(N908),  .B(N940),  .C(add_0_root_add_317_4_carry[6]), .YC(add_0_root_add_317_4_carry[7]), .YS(t1[6]));
   FAX1 add_0_root_add_317_4_U1_7 ( .A(N909),  .B(N941),  .C(add_0_root_add_317_4_carry[7]), .YC(add_0_root_add_317_4_carry[8]), .YS(t1[7]));
   FAX1 add_0_root_add_317_4_U1_8 ( .A(N910),  .B(N942),  .C(add_0_root_add_317_4_carry[8]), .YC(add_0_root_add_317_4_carry[9]), .YS(t1[8]));
   FAX1 add_0_root_add_317_4_U1_9 ( .A(N911),  .B(N943),  .C(add_0_root_add_317_4_carry[9]), .YC(add_0_root_add_317_4_carry[10]), .YS(t1[9]));
   FAX1 add_0_root_add_317_4_U1_10 ( .A(N912),  .B(N944),  .C(add_0_root_add_317_4_carry[10]), .YC(add_0_root_add_317_4_carry[11]), .YS(t1[10]));
   FAX1 add_0_root_add_317_4_U1_11 ( .A(N913),  .B(N945),  .C(add_0_root_add_317_4_carry[11]), .YC(add_0_root_add_317_4_carry[12]), .YS(t1[11]));
   FAX1 add_0_root_add_317_4_U1_12 ( .A(N914),  .B(N946),  .C(add_0_root_add_317_4_carry[12]), .YC(add_0_root_add_317_4_carry[13]), .YS(t1[12]));
   FAX1 add_0_root_add_317_4_U1_13 ( .A(N915),  .B(N947),  .C(add_0_root_add_317_4_carry[13]), .YC(add_0_root_add_317_4_carry[14]), .YS(t1[13]));
   FAX1 add_0_root_add_317_4_U1_14 ( .A(N916),  .B(N948),  .C(add_0_root_add_317_4_carry[14]), .YC(add_0_root_add_317_4_carry[15]), .YS(t1[14]));
   FAX1 add_0_root_add_317_4_U1_15 ( .A(N917),  .B(N949),  .C(add_0_root_add_317_4_carry[15]), .YC(add_0_root_add_317_4_carry[16]), .YS(t1[15]));
   FAX1 add_0_root_add_317_4_U1_16 ( .A(N918),  .B(N950),  .C(add_0_root_add_317_4_carry[16]), .YC(add_0_root_add_317_4_carry[17]), .YS(t1[16]));
   FAX1 add_0_root_add_317_4_U1_17 ( .A(N919),  .B(N951),  .C(add_0_root_add_317_4_carry[17]), .YC(add_0_root_add_317_4_carry[18]), .YS(t1[17]));
   FAX1 add_0_root_add_317_4_U1_18 ( .A(N920),  .B(N952),  .C(add_0_root_add_317_4_carry[18]), .YC(add_0_root_add_317_4_carry[19]), .YS(t1[18]));
   FAX1 add_0_root_add_317_4_U1_19 ( .A(N921),  .B(N953),  .C(add_0_root_add_317_4_carry[19]), .YC(add_0_root_add_317_4_carry[20]), .YS(t1[19]));
   FAX1 add_0_root_add_317_4_U1_20 ( .A(N922),  .B(N954),  .C(add_0_root_add_317_4_carry[20]), .YC(add_0_root_add_317_4_carry[21]), .YS(t1[20]));
   FAX1 add_0_root_add_317_4_U1_21 ( .A(N923),  .B(N955),  .C(add_0_root_add_317_4_carry[21]), .YC(add_0_root_add_317_4_carry[22]), .YS(t1[21]));
   FAX1 add_0_root_add_317_4_U1_22 ( .A(N924),  .B(N956),  .C(add_0_root_add_317_4_carry[22]), .YC(add_0_root_add_317_4_carry[23]), .YS(t1[22]));
   FAX1 add_0_root_add_317_4_U1_23 ( .A(N925),  .B(N957),  .C(add_0_root_add_317_4_carry[23]), .YC(add_0_root_add_317_4_carry[24]), .YS(t1[23]));
   FAX1 add_0_root_add_317_4_U1_24 ( .A(N926),  .B(N958),  .C(add_0_root_add_317_4_carry[24]), .YC(add_0_root_add_317_4_carry[25]), .YS(t1[24]));
   FAX1 add_0_root_add_317_4_U1_25 ( .A(N927),  .B(N959),  .C(add_0_root_add_317_4_carry[25]), .YC(add_0_root_add_317_4_carry[26]), .YS(t1[25]));
   FAX1 add_0_root_add_317_4_U1_26 ( .A(N928),  .B(N960),  .C(add_0_root_add_317_4_carry[26]), .YC(add_0_root_add_317_4_carry[27]), .YS(t1[26]));
   FAX1 add_0_root_add_317_4_U1_27 ( .A(N929),  .B(N961),  .C(add_0_root_add_317_4_carry[27]), .YC(add_0_root_add_317_4_carry[28]), .YS(t1[27]));
   FAX1 add_0_root_add_317_4_U1_28 ( .A(N930),  .B(N962),  .C(add_0_root_add_317_4_carry[28]), .YC(add_0_root_add_317_4_carry[29]), .YS(t1[28]));
   FAX1 add_0_root_add_317_4_U1_29 ( .A(N931),  .B(N963),  .C(add_0_root_add_317_4_carry[29]), .YC(add_0_root_add_317_4_carry[30]), .YS(t1[29]));
   FAX1 add_0_root_add_317_4_U1_30 ( .A(N932),  .B(N964),  .C(add_0_root_add_317_4_carry[30]), .YC(add_0_root_add_317_4_carry[31]), .YS(t1[30]));
   FAX1 add_0_root_add_317_4_U1_31 ( .A(N933),  .B(N965),  .C(add_0_root_add_317_4_carry[31]), .YS(t1[31]));
   FAX1 add_1_root_add_317_4_U1_1 ( .A(n1818),  .B(N871),  .C(n2961), .YC(add_1_root_add_317_4_carry[2]), .YS(N935));
   FAX1 add_1_root_add_317_4_U1_2 ( .A(n1774),  .B(N872),  .C(add_1_root_add_317_4_carry[2]), .YC(add_1_root_add_317_4_carry[3]), .YS(N936));
   FAX1 add_1_root_add_317_4_U1_3 ( .A(n1773),  .B(N873),  .C(add_1_root_add_317_4_carry[3]), .YC(add_1_root_add_317_4_carry[4]), .YS(N937));
   FAX1 add_1_root_add_317_4_U1_4 ( .A(n1772),  .B(N874),  .C(add_1_root_add_317_4_carry[4]), .YC(add_1_root_add_317_4_carry[5]), .YS(N938));
   FAX1 add_1_root_add_317_4_U1_5 ( .A(n1771),  .B(N875),  .C(add_1_root_add_317_4_carry[5]), .YC(add_1_root_add_317_4_carry[6]), .YS(N939));
   FAX1 add_1_root_add_317_4_U1_6 ( .A(k_data[6]),  .B(N876),  .C(add_1_root_add_317_4_carry[6]), .YC(add_1_root_add_317_4_carry[7]), .YS(N940));
   FAX1 add_1_root_add_317_4_U1_7 ( .A(k_data[7]),  .B(N877),  .C(add_1_root_add_317_4_carry[7]), .YC(add_1_root_add_317_4_carry[8]), .YS(N941));
   FAX1 add_1_root_add_317_4_U1_8 ( .A(n1770),  .B(N878),  .C(add_1_root_add_317_4_carry[8]), .YC(add_1_root_add_317_4_carry[9]), .YS(N942));
   FAX1 add_1_root_add_317_4_U1_9 ( .A(n1769),  .B(N879),  .C(add_1_root_add_317_4_carry[9]), .YC(add_1_root_add_317_4_carry[10]), .YS(N943));
   FAX1 add_1_root_add_317_4_U1_10 ( .A(n1768),  .B(N880),  .C(add_1_root_add_317_4_carry[10]), .YC(add_1_root_add_317_4_carry[11]), .YS(N944));
   FAX1 add_1_root_add_317_4_U1_11 ( .A(n2779),  .B(N881),  .C(add_1_root_add_317_4_carry[11]), .YC(add_1_root_add_317_4_carry[12]), .YS(N945));
   FAX1 add_1_root_add_317_4_U1_12 ( .A(k_data[12]),  .B(N882),  .C(add_1_root_add_317_4_carry[12]), .YC(add_1_root_add_317_4_carry[13]), .YS(N946));
   FAX1 add_1_root_add_317_4_U1_13 ( .A(n1767),  .B(N883),  .C(add_1_root_add_317_4_carry[13]), .YC(add_1_root_add_317_4_carry[14]), .YS(N947));
   FAX1 add_1_root_add_317_4_U1_14 ( .A(n1817),  .B(N884),  .C(add_1_root_add_317_4_carry[14]), .YC(add_1_root_add_317_4_carry[15]), .YS(N948));
   FAX1 add_1_root_add_317_4_U1_15 ( .A(n2086),  .B(N885),  .C(add_1_root_add_317_4_carry[15]), .YC(add_1_root_add_317_4_carry[16]), .YS(N949));
   FAX1 add_1_root_add_317_4_U1_16 ( .A(n1766),  .B(N886),  .C(add_1_root_add_317_4_carry[16]), .YC(add_1_root_add_317_4_carry[17]), .YS(N950));
   FAX1 add_1_root_add_317_4_U1_17 ( .A(k_data[17]),  .B(N887),  .C(add_1_root_add_317_4_carry[17]), .YC(add_1_root_add_317_4_carry[18]), .YS(N951));
   FAX1 add_1_root_add_317_4_U1_18 ( .A(n1765),  .B(N888),  .C(add_1_root_add_317_4_carry[18]), .YC(add_1_root_add_317_4_carry[19]), .YS(N952));
   FAX1 add_1_root_add_317_4_U1_19 ( .A(k_data[19]),  .B(N889),  .C(add_1_root_add_317_4_carry[19]), .YC(add_1_root_add_317_4_carry[20]), .YS(N953));
   FAX1 add_1_root_add_317_4_U1_20 ( .A(n2649),  .B(N890),  .C(add_1_root_add_317_4_carry[20]), .YC(add_1_root_add_317_4_carry[21]), .YS(N954));
   FAX1 add_1_root_add_317_4_U1_21 ( .A(n1764),  .B(N891),  .C(add_1_root_add_317_4_carry[21]), .YC(add_1_root_add_317_4_carry[22]), .YS(N955));
   FAX1 add_1_root_add_317_4_U1_22 ( .A(n1763),  .B(N892),  .C(add_1_root_add_317_4_carry[22]), .YC(add_1_root_add_317_4_carry[23]), .YS(N956));
   FAX1 add_1_root_add_317_4_U1_23 ( .A(n2072),  .B(N893),  .C(add_1_root_add_317_4_carry[23]), .YC(add_1_root_add_317_4_carry[24]), .YS(N957));
   FAX1 add_1_root_add_317_4_U1_24 ( .A(n1762),  .B(N894),  .C(add_1_root_add_317_4_carry[24]), .YC(add_1_root_add_317_4_carry[25]), .YS(N958));
   FAX1 add_1_root_add_317_4_U1_25 ( .A(n2537),  .B(N895),  .C(add_1_root_add_317_4_carry[25]), .YC(add_1_root_add_317_4_carry[26]), .YS(N959));
   FAX1 add_1_root_add_317_4_U1_26 ( .A(n2480),  .B(N896),  .C(add_1_root_add_317_4_carry[26]), .YC(add_1_root_add_317_4_carry[27]), .YS(N960));
   FAX1 add_1_root_add_317_4_U1_27 ( .A(n1761),  .B(N897),  .C(add_1_root_add_317_4_carry[27]), .YC(add_1_root_add_317_4_carry[28]), .YS(N961));
   FAX1 add_1_root_add_317_4_U1_28 ( .A(n1760),  .B(N898),  .C(add_1_root_add_317_4_carry[28]), .YC(add_1_root_add_317_4_carry[29]), .YS(N962));
   FAX1 add_1_root_add_317_4_U1_29 ( .A(k_data[29]),  .B(N899),  .C(add_1_root_add_317_4_carry[29]), .YC(add_1_root_add_317_4_carry[30]), .YS(N963));
   FAX1 add_1_root_add_317_4_U1_30 ( .A(k_data[30]),  .B(N900),  .C(add_1_root_add_317_4_carry[30]), .YC(add_1_root_add_317_4_carry[31]), .YS(N964));
   FAX1 add_1_root_add_317_4_U1_31 ( .A(n1816),  .B(N901),  .C(add_1_root_add_317_4_carry[31]), .YS(N965));
   FAX1 add_2_root_add_317_4_U1_1 ( .A(N868),  .B(n1757),  .C(n1850), .YC(add_2_root_add_317_4_carry[2]), .YS(N903));
   FAX1 add_2_root_add_317_4_U1_2 ( .A(N867),  .B(n1848),  .C(add_2_root_add_317_4_carry[2]), .YC(add_2_root_add_317_4_carry[3]), .YS(N904));
   FAX1 add_2_root_add_317_4_U1_3 ( .A(N866),  .B(n1847),  .C(add_2_root_add_317_4_carry[3]), .YC(add_2_root_add_317_4_carry[4]), .YS(N905));
   FAX1 add_2_root_add_317_4_U1_4 ( .A(N865),  .B(n1846),  .C(add_2_root_add_317_4_carry[4]), .YC(add_2_root_add_317_4_carry[5]), .YS(N906));
   FAX1 add_2_root_add_317_4_U1_5 ( .A(N864),  .B(n1845),  .C(add_2_root_add_317_4_carry[5]), .YC(add_2_root_add_317_4_carry[6]), .YS(N907));
   FAX1 add_2_root_add_317_4_U1_6 ( .A(N863),  .B(n1844),  .C(add_2_root_add_317_4_carry[6]), .YC(add_2_root_add_317_4_carry[7]), .YS(N908));
   FAX1 add_2_root_add_317_4_U1_7 ( .A(N862),  .B(n1843),  .C(add_2_root_add_317_4_carry[7]), .YC(add_2_root_add_317_4_carry[8]), .YS(N909));
   FAX1 add_2_root_add_317_4_U1_8 ( .A(N861),  .B(n1842),  .C(add_2_root_add_317_4_carry[8]), .YC(add_2_root_add_317_4_carry[9]), .YS(N910));
   FAX1 add_2_root_add_317_4_U1_9 ( .A(N860),  .B(n1841),  .C(add_2_root_add_317_4_carry[9]), .YC(add_2_root_add_317_4_carry[10]), .YS(N911));
   FAX1 add_2_root_add_317_4_U1_10 ( .A(N859),  .B(n1830),  .C(add_2_root_add_317_4_carry[10]), .YC(add_2_root_add_317_4_carry[11]), .YS(N912));
   FAX1 add_2_root_add_317_4_U1_11 ( .A(N858),  .B(n1829),  .C(add_2_root_add_317_4_carry[11]), .YC(add_2_root_add_317_4_carry[12]), .YS(N913));
   FAX1 add_2_root_add_317_4_U1_12 ( .A(N857),  .B(n1828),  .C(add_2_root_add_317_4_carry[12]), .YC(add_2_root_add_317_4_carry[13]), .YS(N914));
   FAX1 add_2_root_add_317_4_U1_13 ( .A(N856),  .B(n1827),  .C(add_2_root_add_317_4_carry[13]), .YC(add_2_root_add_317_4_carry[14]), .YS(N915));
   FAX1 add_2_root_add_317_4_U1_14 ( .A(N855),  .B(n1826),  .C(add_2_root_add_317_4_carry[14]), .YC(add_2_root_add_317_4_carry[15]), .YS(N916));
   FAX1 add_2_root_add_317_4_U1_15 ( .A(N854),  .B(n1825),  .C(add_2_root_add_317_4_carry[15]), .YC(add_2_root_add_317_4_carry[16]), .YS(N917));
   FAX1 add_2_root_add_317_4_U1_16 ( .A(N853),  .B(n1824),  .C(add_2_root_add_317_4_carry[16]), .YC(add_2_root_add_317_4_carry[17]), .YS(N918));
   FAX1 add_2_root_add_317_4_U1_17 ( .A(N852),  .B(n1823),  .C(add_2_root_add_317_4_carry[17]), .YC(add_2_root_add_317_4_carry[18]), .YS(N919));
   FAX1 add_2_root_add_317_4_U1_18 ( .A(N851),  .B(n1822),  .C(add_2_root_add_317_4_carry[18]), .YC(add_2_root_add_317_4_carry[19]), .YS(N920));
   FAX1 add_2_root_add_317_4_U1_19 ( .A(N850),  .B(n1821),  .C(add_2_root_add_317_4_carry[19]), .YC(add_2_root_add_317_4_carry[20]), .YS(N921));
   FAX1 add_2_root_add_317_4_U1_20 ( .A(N849),  .B(n1820),  .C(add_2_root_add_317_4_carry[20]), .YC(add_2_root_add_317_4_carry[21]), .YS(N922));
   FAX1 add_2_root_add_317_4_U1_21 ( .A(N848),  .B(n1819),  .C(add_2_root_add_317_4_carry[21]), .YC(add_2_root_add_317_4_carry[22]), .YS(N923));
   FAX1 add_2_root_add_317_4_U1_22 ( .A(N847),  .B(n1840),  .C(add_2_root_add_317_4_carry[22]), .YC(add_2_root_add_317_4_carry[23]), .YS(N924));
   FAX1 add_2_root_add_317_4_U1_23 ( .A(N846),  .B(n1839),  .C(add_2_root_add_317_4_carry[23]), .YC(add_2_root_add_317_4_carry[24]), .YS(N925));
   FAX1 add_2_root_add_317_4_U1_24 ( .A(N845),  .B(n1838),  .C(add_2_root_add_317_4_carry[24]), .YC(add_2_root_add_317_4_carry[25]), .YS(N926));
   FAX1 add_2_root_add_317_4_U1_25 ( .A(N844),  .B(n1837),  .C(add_2_root_add_317_4_carry[25]), .YC(add_2_root_add_317_4_carry[26]), .YS(N927));
   FAX1 add_2_root_add_317_4_U1_26 ( .A(N843),  .B(n1836),  .C(add_2_root_add_317_4_carry[26]), .YC(add_2_root_add_317_4_carry[27]), .YS(N928));
   FAX1 add_2_root_add_317_4_U1_27 ( .A(N842),  .B(n1835),  .C(add_2_root_add_317_4_carry[27]), .YC(add_2_root_add_317_4_carry[28]), .YS(N929));
   FAX1 add_2_root_add_317_4_U1_28 ( .A(N841),  .B(n1834),  .C(add_2_root_add_317_4_carry[28]), .YC(add_2_root_add_317_4_carry[29]), .YS(N930));
   FAX1 add_2_root_add_317_4_U1_29 ( .A(N840),  .B(n1833),  .C(add_2_root_add_317_4_carry[29]), .YC(add_2_root_add_317_4_carry[30]), .YS(N931));
   FAX1 add_2_root_add_317_4_U1_30 ( .A(N839),  .B(n1832),  .C(add_2_root_add_317_4_carry[30]), .YC(add_2_root_add_317_4_carry[31]), .YS(N932));
   FAX1 add_2_root_add_317_4_U1_31 ( .A(N838),  .B(n1831),  .C(add_2_root_add_317_4_carry[31]), .YS(N933));
   FAX1 add_3_root_add_317_4_U1_1 ( .A(h_reg[1]),  .B(N836),  .C(n2966), .YC(add_3_root_add_317_4_carry[2]), .YS(N871));
   FAX1 add_3_root_add_317_4_U1_2 ( .A(h_reg[2]),  .B(N835),  .C(add_3_root_add_317_4_carry[2]), .YC(add_3_root_add_317_4_carry[3]), .YS(N872));
   FAX1 add_3_root_add_317_4_U1_3 ( .A(h_reg[3]),  .B(N834),  .C(add_3_root_add_317_4_carry[3]), .YC(add_3_root_add_317_4_carry[4]), .YS(N873));
   FAX1 add_3_root_add_317_4_U1_4 ( .A(h_reg[4]),  .B(N833),  .C(add_3_root_add_317_4_carry[4]), .YC(add_3_root_add_317_4_carry[5]), .YS(N874));
   FAX1 add_3_root_add_317_4_U1_5 ( .A(h_reg[5]),  .B(N832),  .C(add_3_root_add_317_4_carry[5]), .YC(add_3_root_add_317_4_carry[6]), .YS(N875));
   FAX1 add_3_root_add_317_4_U1_6 ( .A(h_reg[6]),  .B(N831),  .C(add_3_root_add_317_4_carry[6]), .YC(add_3_root_add_317_4_carry[7]), .YS(N876));
   FAX1 add_3_root_add_317_4_U1_7 ( .A(h_reg[7]),  .B(N830),  .C(add_3_root_add_317_4_carry[7]), .YC(add_3_root_add_317_4_carry[8]), .YS(N877));
   FAX1 add_3_root_add_317_4_U1_8 ( .A(h_reg[8]),  .B(N829),  .C(add_3_root_add_317_4_carry[8]), .YC(add_3_root_add_317_4_carry[9]), .YS(N878));
   FAX1 add_3_root_add_317_4_U1_9 ( .A(h_reg[9]),  .B(N828),  .C(add_3_root_add_317_4_carry[9]), .YC(add_3_root_add_317_4_carry[10]), .YS(N879));
   FAX1 add_3_root_add_317_4_U1_10 ( .A(h_reg[10]),  .B(N827),  .C(add_3_root_add_317_4_carry[10]), .YC(add_3_root_add_317_4_carry[11]), .YS(N880));
   FAX1 add_3_root_add_317_4_U1_11 ( .A(h_reg[11]),  .B(N826),  .C(add_3_root_add_317_4_carry[11]), .YC(add_3_root_add_317_4_carry[12]), .YS(N881));
   FAX1 add_3_root_add_317_4_U1_12 ( .A(h_reg[12]),  .B(N825),  .C(add_3_root_add_317_4_carry[12]), .YC(add_3_root_add_317_4_carry[13]), .YS(N882));
   FAX1 add_3_root_add_317_4_U1_13 ( .A(h_reg[13]),  .B(N824),  .C(add_3_root_add_317_4_carry[13]), .YC(add_3_root_add_317_4_carry[14]), .YS(N883));
   FAX1 add_3_root_add_317_4_U1_14 ( .A(h_reg[14]),  .B(N823),  .C(add_3_root_add_317_4_carry[14]), .YC(add_3_root_add_317_4_carry[15]), .YS(N884));
   FAX1 add_3_root_add_317_4_U1_15 ( .A(h_reg[15]),  .B(N822),  .C(add_3_root_add_317_4_carry[15]), .YC(add_3_root_add_317_4_carry[16]), .YS(N885));
   FAX1 add_3_root_add_317_4_U1_16 ( .A(h_reg[16]),  .B(N821),  .C(add_3_root_add_317_4_carry[16]), .YC(add_3_root_add_317_4_carry[17]), .YS(N886));
   FAX1 add_3_root_add_317_4_U1_17 ( .A(h_reg[17]),  .B(N820),  .C(add_3_root_add_317_4_carry[17]), .YC(add_3_root_add_317_4_carry[18]), .YS(N887));
   FAX1 add_3_root_add_317_4_U1_18 ( .A(h_reg[18]),  .B(N819),  .C(add_3_root_add_317_4_carry[18]), .YC(add_3_root_add_317_4_carry[19]), .YS(N888));
   FAX1 add_3_root_add_317_4_U1_19 ( .A(h_reg[19]),  .B(N818),  .C(add_3_root_add_317_4_carry[19]), .YC(add_3_root_add_317_4_carry[20]), .YS(N889));
   FAX1 add_3_root_add_317_4_U1_20 ( .A(h_reg[20]),  .B(N817),  .C(add_3_root_add_317_4_carry[20]), .YC(add_3_root_add_317_4_carry[21]), .YS(N890));
   FAX1 add_3_root_add_317_4_U1_21 ( .A(h_reg[21]),  .B(N816),  .C(add_3_root_add_317_4_carry[21]), .YC(add_3_root_add_317_4_carry[22]), .YS(N891));
   FAX1 add_3_root_add_317_4_U1_22 ( .A(h_reg[22]),  .B(N815),  .C(add_3_root_add_317_4_carry[22]), .YC(add_3_root_add_317_4_carry[23]), .YS(N892));
   FAX1 add_3_root_add_317_4_U1_23 ( .A(h_reg[23]),  .B(N814),  .C(add_3_root_add_317_4_carry[23]), .YC(add_3_root_add_317_4_carry[24]), .YS(N893));
   FAX1 add_3_root_add_317_4_U1_24 ( .A(h_reg[24]),  .B(N813),  .C(add_3_root_add_317_4_carry[24]), .YC(add_3_root_add_317_4_carry[25]), .YS(N894));
   FAX1 add_3_root_add_317_4_U1_25 ( .A(h_reg[25]),  .B(N812),  .C(add_3_root_add_317_4_carry[25]), .YC(add_3_root_add_317_4_carry[26]), .YS(N895));
   FAX1 add_3_root_add_317_4_U1_26 ( .A(h_reg[26]),  .B(N811),  .C(add_3_root_add_317_4_carry[26]), .YC(add_3_root_add_317_4_carry[27]), .YS(N896));
   FAX1 add_3_root_add_317_4_U1_27 ( .A(h_reg[27]),  .B(N810),  .C(add_3_root_add_317_4_carry[27]), .YC(add_3_root_add_317_4_carry[28]), .YS(N897));
   FAX1 add_3_root_add_317_4_U1_28 ( .A(h_reg[28]),  .B(N809),  .C(add_3_root_add_317_4_carry[28]), .YC(add_3_root_add_317_4_carry[29]), .YS(N898));
   FAX1 add_3_root_add_317_4_U1_29 ( .A(h_reg[29]),  .B(N808),  .C(add_3_root_add_317_4_carry[29]), .YC(add_3_root_add_317_4_carry[30]), .YS(N899));
   FAX1 add_3_root_add_317_4_U1_30 ( .A(h_reg[30]),  .B(N807),  .C(add_3_root_add_317_4_carry[30]), .YC(add_3_root_add_317_4_carry[31]), .YS(N900));
   FAX1 add_3_root_add_317_4_U1_31 ( .A(h_reg[31]),  .B(N806),  .C(add_3_root_add_317_4_carry[31]), .YS(N901));
   FAX1 add_295_U1_1 ( .A(digest[1]),  .B(h_reg[1]),  .C(n2969), .YC(add_295_carry[2]), .YS(N775));
   FAX1 add_295_U1_2 ( .A(digest[2]),  .B(h_reg[2]),  .C(add_295_carry[2]), .YC(add_295_carry[3]), .YS(N776));
   FAX1 add_295_U1_3 ( .A(digest[3]),  .B(h_reg[3]),  .C(add_295_carry[3]), .YC(add_295_carry[4]), .YS(N777));
   FAX1 add_295_U1_4 ( .A(digest[4]),  .B(h_reg[4]),  .C(add_295_carry[4]), .YC(add_295_carry[5]), .YS(N778));
   FAX1 add_295_U1_5 ( .A(digest[5]),  .B(h_reg[5]),  .C(add_295_carry[5]), .YC(add_295_carry[6]), .YS(N779));
   FAX1 add_295_U1_6 ( .A(digest[6]),  .B(h_reg[6]),  .C(add_295_carry[6]), .YC(add_295_carry[7]), .YS(N780));
   FAX1 add_295_U1_7 ( .A(digest[7]),  .B(h_reg[7]),  .C(add_295_carry[7]), .YC(add_295_carry[8]), .YS(N781));
   FAX1 add_295_U1_8 ( .A(digest[8]),  .B(h_reg[8]),  .C(add_295_carry[8]), .YC(add_295_carry[9]), .YS(N782));
   FAX1 add_295_U1_9 ( .A(digest[9]),  .B(h_reg[9]),  .C(add_295_carry[9]), .YC(add_295_carry[10]), .YS(N783));
   FAX1 add_295_U1_10 ( .A(digest[10]),  .B(h_reg[10]),  .C(add_295_carry[10]), .YC(add_295_carry[11]), .YS(N784));
   FAX1 add_295_U1_11 ( .A(digest[11]),  .B(h_reg[11]),  .C(add_295_carry[11]), .YC(add_295_carry[12]), .YS(N785));
   FAX1 add_295_U1_12 ( .A(digest[12]),  .B(h_reg[12]),  .C(add_295_carry[12]), .YC(add_295_carry[13]), .YS(N786));
   FAX1 add_295_U1_13 ( .A(digest[13]),  .B(h_reg[13]),  .C(add_295_carry[13]), .YC(add_295_carry[14]), .YS(N787));
   FAX1 add_295_U1_14 ( .A(digest[14]),  .B(h_reg[14]),  .C(add_295_carry[14]), .YC(add_295_carry[15]), .YS(N788));
   FAX1 add_295_U1_15 ( .A(digest[15]),  .B(h_reg[15]),  .C(add_295_carry[15]), .YC(add_295_carry[16]), .YS(N789));
   FAX1 add_295_U1_16 ( .A(digest[16]),  .B(h_reg[16]),  .C(add_295_carry[16]), .YC(add_295_carry[17]), .YS(N790));
   FAX1 add_295_U1_17 ( .A(digest[17]),  .B(h_reg[17]),  .C(add_295_carry[17]), .YC(add_295_carry[18]), .YS(N791));
   FAX1 add_295_U1_18 ( .A(digest[18]),  .B(h_reg[18]),  .C(add_295_carry[18]), .YC(add_295_carry[19]), .YS(N792));
   FAX1 add_295_U1_19 ( .A(digest[19]),  .B(h_reg[19]),  .C(add_295_carry[19]), .YC(add_295_carry[20]), .YS(N793));
   FAX1 add_295_U1_20 ( .A(digest[20]),  .B(h_reg[20]),  .C(add_295_carry[20]), .YC(add_295_carry[21]), .YS(N794));
   FAX1 add_295_U1_21 ( .A(digest[21]),  .B(h_reg[21]),  .C(add_295_carry[21]), .YC(add_295_carry[22]), .YS(N795));
   FAX1 add_295_U1_22 ( .A(digest[22]),  .B(h_reg[22]),  .C(add_295_carry[22]), .YC(add_295_carry[23]), .YS(N796));
   FAX1 add_295_U1_23 ( .A(digest[23]),  .B(h_reg[23]),  .C(add_295_carry[23]), .YC(add_295_carry[24]), .YS(N797));
   FAX1 add_295_U1_24 ( .A(digest[24]),  .B(h_reg[24]),  .C(add_295_carry[24]), .YC(add_295_carry[25]), .YS(N798));
   FAX1 add_295_U1_25 ( .A(digest[25]),  .B(h_reg[25]),  .C(add_295_carry[25]), .YC(add_295_carry[26]), .YS(N799));
   FAX1 add_295_U1_26 ( .A(digest[26]),  .B(h_reg[26]),  .C(add_295_carry[26]), .YC(add_295_carry[27]), .YS(N800));
   FAX1 add_295_U1_27 ( .A(digest[27]),  .B(h_reg[27]),  .C(add_295_carry[27]), .YC(add_295_carry[28]), .YS(N801));
   FAX1 add_295_U1_28 ( .A(digest[28]),  .B(h_reg[28]),  .C(add_295_carry[28]), .YC(add_295_carry[29]), .YS(N802));
   FAX1 add_295_U1_29 ( .A(digest[29]),  .B(h_reg[29]),  .C(add_295_carry[29]), .YC(add_295_carry[30]), .YS(N803));
   FAX1 add_295_U1_30 ( .A(digest[30]),  .B(h_reg[30]),  .C(add_295_carry[30]), .YC(add_295_carry[31]), .YS(N804));
   FAX1 add_295_U1_31 ( .A(digest[31]),  .B(h_reg[31]),  .C(add_295_carry[31]), .YS(N805));
   FAX1 add_294_U1_1 ( .A(digest[33]),  .B(g_reg[1]),  .C(n2974), .YC(add_294_carry[2]), .YS(N743));
   FAX1 add_294_U1_2 ( .A(digest[34]),  .B(g_reg[2]),  .C(add_294_carry[2]), .YC(add_294_carry[3]), .YS(N744));
   FAX1 add_294_U1_3 ( .A(digest[35]),  .B(g_reg[3]),  .C(add_294_carry[3]), .YC(add_294_carry[4]), .YS(N745));
   FAX1 add_294_U1_4 ( .A(digest[36]),  .B(g_reg[4]),  .C(add_294_carry[4]), .YC(add_294_carry[5]), .YS(N746));
   FAX1 add_294_U1_5 ( .A(digest[37]),  .B(g_reg[5]),  .C(add_294_carry[5]), .YC(add_294_carry[6]), .YS(N747));
   FAX1 add_294_U1_6 ( .A(digest[38]),  .B(g_reg[6]),  .C(add_294_carry[6]), .YC(add_294_carry[7]), .YS(N748));
   FAX1 add_294_U1_7 ( .A(digest[39]),  .B(g_reg[7]),  .C(add_294_carry[7]), .YC(add_294_carry[8]), .YS(N749));
   FAX1 add_294_U1_8 ( .A(digest[40]),  .B(g_reg[8]),  .C(add_294_carry[8]), .YC(add_294_carry[9]), .YS(N750));
   FAX1 add_294_U1_9 ( .A(digest[41]),  .B(g_reg[9]),  .C(add_294_carry[9]), .YC(add_294_carry[10]), .YS(N751));
   FAX1 add_294_U1_10 ( .A(digest[42]),  .B(g_reg[10]),  .C(add_294_carry[10]), .YC(add_294_carry[11]), .YS(N752));
   FAX1 add_294_U1_11 ( .A(digest[43]),  .B(g_reg[11]),  .C(add_294_carry[11]), .YC(add_294_carry[12]), .YS(N753));
   FAX1 add_294_U1_12 ( .A(digest[44]),  .B(g_reg[12]),  .C(add_294_carry[12]), .YC(add_294_carry[13]), .YS(N754));
   FAX1 add_294_U1_13 ( .A(digest[45]),  .B(g_reg[13]),  .C(add_294_carry[13]), .YC(add_294_carry[14]), .YS(N755));
   FAX1 add_294_U1_14 ( .A(digest[46]),  .B(g_reg[14]),  .C(add_294_carry[14]), .YC(add_294_carry[15]), .YS(N756));
   FAX1 add_294_U1_15 ( .A(digest[47]),  .B(g_reg[15]),  .C(add_294_carry[15]), .YC(add_294_carry[16]), .YS(N757));
   FAX1 add_294_U1_16 ( .A(digest[48]),  .B(g_reg[16]),  .C(add_294_carry[16]), .YC(add_294_carry[17]), .YS(N758));
   FAX1 add_294_U1_17 ( .A(digest[49]),  .B(g_reg[17]),  .C(add_294_carry[17]), .YC(add_294_carry[18]), .YS(N759));
   FAX1 add_294_U1_18 ( .A(digest[50]),  .B(g_reg[18]),  .C(add_294_carry[18]), .YC(add_294_carry[19]), .YS(N760));
   FAX1 add_294_U1_19 ( .A(digest[51]),  .B(g_reg[19]),  .C(add_294_carry[19]), .YC(add_294_carry[20]), .YS(N761));
   FAX1 add_294_U1_20 ( .A(digest[52]),  .B(g_reg[20]),  .C(add_294_carry[20]), .YC(add_294_carry[21]), .YS(N762));
   FAX1 add_294_U1_21 ( .A(digest[53]),  .B(g_reg[21]),  .C(add_294_carry[21]), .YC(add_294_carry[22]), .YS(N763));
   FAX1 add_294_U1_22 ( .A(digest[54]),  .B(g_reg[22]),  .C(add_294_carry[22]), .YC(add_294_carry[23]), .YS(N764));
   FAX1 add_294_U1_23 ( .A(digest[55]),  .B(g_reg[23]),  .C(add_294_carry[23]), .YC(add_294_carry[24]), .YS(N765));
   FAX1 add_294_U1_24 ( .A(digest[56]),  .B(g_reg[24]),  .C(add_294_carry[24]), .YC(add_294_carry[25]), .YS(N766));
   FAX1 add_294_U1_25 ( .A(digest[57]),  .B(g_reg[25]),  .C(add_294_carry[25]), .YC(add_294_carry[26]), .YS(N767));
   FAX1 add_294_U1_26 ( .A(digest[58]),  .B(g_reg[26]),  .C(add_294_carry[26]), .YC(add_294_carry[27]), .YS(N768));
   FAX1 add_294_U1_27 ( .A(digest[59]),  .B(g_reg[27]),  .C(add_294_carry[27]), .YC(add_294_carry[28]), .YS(N769));
   FAX1 add_294_U1_28 ( .A(digest[60]),  .B(g_reg[28]),  .C(add_294_carry[28]), .YC(add_294_carry[29]), .YS(N770));
   FAX1 add_294_U1_29 ( .A(digest[61]),  .B(g_reg[29]),  .C(add_294_carry[29]), .YC(add_294_carry[30]), .YS(N771));
   FAX1 add_294_U1_30 ( .A(digest[62]),  .B(g_reg[30]),  .C(add_294_carry[30]), .YC(add_294_carry[31]), .YS(N772));
   FAX1 add_294_U1_31 ( .A(digest[63]),  .B(g_reg[31]),  .C(add_294_carry[31]), .YS(N773));
   FAX1 add_293_U1_1 ( .A(digest[65]),  .B(f_reg[1]),  .C(n2970), .YC(add_293_carry[2]), .YS(N711));
   FAX1 add_293_U1_2 ( .A(digest[66]),  .B(f_reg[2]),  .C(add_293_carry[2]), .YC(add_293_carry[3]), .YS(N712));
   FAX1 add_293_U1_3 ( .A(digest[67]),  .B(f_reg[3]),  .C(add_293_carry[3]), .YC(add_293_carry[4]), .YS(N713));
   FAX1 add_293_U1_4 ( .A(digest[68]),  .B(f_reg[4]),  .C(add_293_carry[4]), .YC(add_293_carry[5]), .YS(N714));
   FAX1 add_293_U1_5 ( .A(digest[69]),  .B(f_reg[5]),  .C(add_293_carry[5]), .YC(add_293_carry[6]), .YS(N715));
   FAX1 add_293_U1_6 ( .A(digest[70]),  .B(f_reg[6]),  .C(add_293_carry[6]), .YC(add_293_carry[7]), .YS(N716));
   FAX1 add_293_U1_7 ( .A(digest[71]),  .B(f_reg[7]),  .C(add_293_carry[7]), .YC(add_293_carry[8]), .YS(N717));
   FAX1 add_293_U1_8 ( .A(digest[72]),  .B(f_reg[8]),  .C(add_293_carry[8]), .YC(add_293_carry[9]), .YS(N718));
   FAX1 add_293_U1_9 ( .A(digest[73]),  .B(f_reg[9]),  .C(add_293_carry[9]), .YC(add_293_carry[10]), .YS(N719));
   FAX1 add_293_U1_10 ( .A(digest[74]),  .B(f_reg[10]),  .C(add_293_carry[10]), .YC(add_293_carry[11]), .YS(N720));
   FAX1 add_293_U1_11 ( .A(digest[75]),  .B(f_reg[11]),  .C(add_293_carry[11]), .YC(add_293_carry[12]), .YS(N721));
   FAX1 add_293_U1_12 ( .A(digest[76]),  .B(f_reg[12]),  .C(add_293_carry[12]), .YC(add_293_carry[13]), .YS(N722));
   FAX1 add_293_U1_13 ( .A(digest[77]),  .B(f_reg[13]),  .C(add_293_carry[13]), .YC(add_293_carry[14]), .YS(N723));
   FAX1 add_293_U1_14 ( .A(digest[78]),  .B(f_reg[14]),  .C(add_293_carry[14]), .YC(add_293_carry[15]), .YS(N724));
   FAX1 add_293_U1_15 ( .A(digest[79]),  .B(f_reg[15]),  .C(add_293_carry[15]), .YC(add_293_carry[16]), .YS(N725));
   FAX1 add_293_U1_16 ( .A(digest[80]),  .B(f_reg[16]),  .C(add_293_carry[16]), .YC(add_293_carry[17]), .YS(N726));
   FAX1 add_293_U1_17 ( .A(digest[81]),  .B(f_reg[17]),  .C(add_293_carry[17]), .YC(add_293_carry[18]), .YS(N727));
   FAX1 add_293_U1_18 ( .A(digest[82]),  .B(f_reg[18]),  .C(add_293_carry[18]), .YC(add_293_carry[19]), .YS(N728));
   FAX1 add_293_U1_19 ( .A(digest[83]),  .B(f_reg[19]),  .C(add_293_carry[19]), .YC(add_293_carry[20]), .YS(N729));
   FAX1 add_293_U1_20 ( .A(digest[84]),  .B(f_reg[20]),  .C(add_293_carry[20]), .YC(add_293_carry[21]), .YS(N730));
   FAX1 add_293_U1_21 ( .A(digest[85]),  .B(f_reg[21]),  .C(add_293_carry[21]), .YC(add_293_carry[22]), .YS(N731));
   FAX1 add_293_U1_22 ( .A(digest[86]),  .B(f_reg[22]),  .C(add_293_carry[22]), .YC(add_293_carry[23]), .YS(N732));
   FAX1 add_293_U1_23 ( .A(digest[87]),  .B(f_reg[23]),  .C(add_293_carry[23]), .YC(add_293_carry[24]), .YS(N733));
   FAX1 add_293_U1_24 ( .A(digest[88]),  .B(f_reg[24]),  .C(add_293_carry[24]), .YC(add_293_carry[25]), .YS(N734));
   FAX1 add_293_U1_25 ( .A(digest[89]),  .B(f_reg[25]),  .C(add_293_carry[25]), .YC(add_293_carry[26]), .YS(N735));
   FAX1 add_293_U1_26 ( .A(digest[90]),  .B(f_reg[26]),  .C(add_293_carry[26]), .YC(add_293_carry[27]), .YS(N736));
   FAX1 add_293_U1_27 ( .A(digest[91]),  .B(f_reg[27]),  .C(add_293_carry[27]), .YC(add_293_carry[28]), .YS(N737));
   FAX1 add_293_U1_28 ( .A(digest[92]),  .B(f_reg[28]),  .C(add_293_carry[28]), .YC(add_293_carry[29]), .YS(N738));
   FAX1 add_293_U1_29 ( .A(digest[93]),  .B(f_reg[29]),  .C(add_293_carry[29]), .YC(add_293_carry[30]), .YS(N739));
   FAX1 add_293_U1_30 ( .A(digest[94]),  .B(f_reg[30]),  .C(add_293_carry[30]), .YC(add_293_carry[31]), .YS(N740));
   FAX1 add_293_U1_31 ( .A(digest[95]),  .B(f_reg[31]),  .C(add_293_carry[31]), .YS(N741));
   FAX1 add_292_U1_1 ( .A(digest[97]),  .B(e_reg[1]),  .C(n2975), .YC(add_292_carry[2]), .YS(N679));
   FAX1 add_292_U1_2 ( .A(digest[98]),  .B(e_reg[2]),  .C(add_292_carry[2]), .YC(add_292_carry[3]), .YS(N680));
   FAX1 add_292_U1_3 ( .A(digest[99]),  .B(e_reg[3]),  .C(add_292_carry[3]), .YC(add_292_carry[4]), .YS(N681));
   FAX1 add_292_U1_4 ( .A(digest[100]),  .B(e_reg[4]),  .C(add_292_carry[4]), .YC(add_292_carry[5]), .YS(N682));
   FAX1 add_292_U1_5 ( .A(digest[101]),  .B(e_reg[5]),  .C(add_292_carry[5]), .YC(add_292_carry[6]), .YS(N683));
   FAX1 add_292_U1_6 ( .A(digest[102]),  .B(e_reg[6]),  .C(add_292_carry[6]), .YC(add_292_carry[7]), .YS(N684));
   FAX1 add_292_U1_7 ( .A(digest[103]),  .B(e_reg[7]),  .C(add_292_carry[7]), .YC(add_292_carry[8]), .YS(N685));
   FAX1 add_292_U1_8 ( .A(digest[104]),  .B(e_reg[8]),  .C(add_292_carry[8]), .YC(add_292_carry[9]), .YS(N686));
   FAX1 add_292_U1_9 ( .A(digest[105]),  .B(e_reg[9]),  .C(add_292_carry[9]), .YC(add_292_carry[10]), .YS(N687));
   FAX1 add_292_U1_10 ( .A(digest[106]),  .B(e_reg[10]),  .C(add_292_carry[10]), .YC(add_292_carry[11]), .YS(N688));
   FAX1 add_292_U1_11 ( .A(digest[107]),  .B(e_reg[11]),  .C(add_292_carry[11]), .YC(add_292_carry[12]), .YS(N689));
   FAX1 add_292_U1_12 ( .A(digest[108]),  .B(e_reg[12]),  .C(add_292_carry[12]), .YC(add_292_carry[13]), .YS(N690));
   FAX1 add_292_U1_13 ( .A(digest[109]),  .B(e_reg[13]),  .C(add_292_carry[13]), .YC(add_292_carry[14]), .YS(N691));
   FAX1 add_292_U1_14 ( .A(digest[110]),  .B(e_reg[14]),  .C(add_292_carry[14]), .YC(add_292_carry[15]), .YS(N692));
   FAX1 add_292_U1_15 ( .A(digest[111]),  .B(e_reg[15]),  .C(add_292_carry[15]), .YC(add_292_carry[16]), .YS(N693));
   FAX1 add_292_U1_16 ( .A(digest[112]),  .B(e_reg[16]),  .C(add_292_carry[16]), .YC(add_292_carry[17]), .YS(N694));
   FAX1 add_292_U1_17 ( .A(digest[113]),  .B(e_reg[17]),  .C(add_292_carry[17]), .YC(add_292_carry[18]), .YS(N695));
   FAX1 add_292_U1_18 ( .A(digest[114]),  .B(e_reg[18]),  .C(add_292_carry[18]), .YC(add_292_carry[19]), .YS(N696));
   FAX1 add_292_U1_19 ( .A(digest[115]),  .B(e_reg[19]),  .C(add_292_carry[19]), .YC(add_292_carry[20]), .YS(N697));
   FAX1 add_292_U1_20 ( .A(digest[116]),  .B(e_reg[20]),  .C(add_292_carry[20]), .YC(add_292_carry[21]), .YS(N698));
   FAX1 add_292_U1_21 ( .A(digest[117]),  .B(e_reg[21]),  .C(add_292_carry[21]), .YC(add_292_carry[22]), .YS(N699));
   FAX1 add_292_U1_22 ( .A(digest[118]),  .B(e_reg[22]),  .C(add_292_carry[22]), .YC(add_292_carry[23]), .YS(N700));
   FAX1 add_292_U1_23 ( .A(digest[119]),  .B(e_reg[23]),  .C(add_292_carry[23]), .YC(add_292_carry[24]), .YS(N701));
   FAX1 add_292_U1_24 ( .A(digest[120]),  .B(e_reg[24]),  .C(add_292_carry[24]), .YC(add_292_carry[25]), .YS(N702));
   FAX1 add_292_U1_25 ( .A(digest[121]),  .B(e_reg[25]),  .C(add_292_carry[25]), .YC(add_292_carry[26]), .YS(N703));
   FAX1 add_292_U1_26 ( .A(digest[122]),  .B(e_reg[26]),  .C(add_292_carry[26]), .YC(add_292_carry[27]), .YS(N704));
   FAX1 add_292_U1_27 ( .A(digest[123]),  .B(e_reg[27]),  .C(add_292_carry[27]), .YC(add_292_carry[28]), .YS(N705));
   FAX1 add_292_U1_28 ( .A(digest[124]),  .B(e_reg[28]),  .C(add_292_carry[28]), .YC(add_292_carry[29]), .YS(N706));
   FAX1 add_292_U1_29 ( .A(digest[125]),  .B(e_reg[29]),  .C(add_292_carry[29]), .YC(add_292_carry[30]), .YS(N707));
   FAX1 add_292_U1_30 ( .A(digest[126]),  .B(e_reg[30]),  .C(add_292_carry[30]), .YC(add_292_carry[31]), .YS(N708));
   FAX1 add_292_U1_31 ( .A(digest[127]),  .B(e_reg[31]),  .C(add_292_carry[31]), .YS(N709));
   FAX1 add_291_U1_1 ( .A(digest[129]),  .B(d_reg[1]),  .C(n2971), .YC(add_291_carry[2]), .YS(N647));
   FAX1 add_291_U1_2 ( .A(digest[130]),  .B(d_reg[2]),  .C(add_291_carry[2]), .YC(add_291_carry[3]), .YS(N648));
   FAX1 add_291_U1_3 ( .A(digest[131]),  .B(d_reg[3]),  .C(add_291_carry[3]), .YC(add_291_carry[4]), .YS(N649));
   FAX1 add_291_U1_4 ( .A(digest[132]),  .B(d_reg[4]),  .C(add_291_carry[4]), .YC(add_291_carry[5]), .YS(N650));
   FAX1 add_291_U1_5 ( .A(digest[133]),  .B(d_reg[5]),  .C(add_291_carry[5]), .YC(add_291_carry[6]), .YS(N651));
   FAX1 add_291_U1_6 ( .A(digest[134]),  .B(d_reg[6]),  .C(add_291_carry[6]), .YC(add_291_carry[7]), .YS(N652));
   FAX1 add_291_U1_7 ( .A(digest[135]),  .B(d_reg[7]),  .C(add_291_carry[7]), .YC(add_291_carry[8]), .YS(N653));
   FAX1 add_291_U1_8 ( .A(digest[136]),  .B(d_reg[8]),  .C(add_291_carry[8]), .YC(add_291_carry[9]), .YS(N654));
   FAX1 add_291_U1_9 ( .A(digest[137]),  .B(d_reg[9]),  .C(add_291_carry[9]), .YC(add_291_carry[10]), .YS(N655));
   FAX1 add_291_U1_10 ( .A(digest[138]),  .B(d_reg[10]),  .C(add_291_carry[10]), .YC(add_291_carry[11]), .YS(N656));
   FAX1 add_291_U1_11 ( .A(digest[139]),  .B(d_reg[11]),  .C(add_291_carry[11]), .YC(add_291_carry[12]), .YS(N657));
   FAX1 add_291_U1_12 ( .A(digest[140]),  .B(d_reg[12]),  .C(add_291_carry[12]), .YC(add_291_carry[13]), .YS(N658));
   FAX1 add_291_U1_13 ( .A(digest[141]),  .B(d_reg[13]),  .C(add_291_carry[13]), .YC(add_291_carry[14]), .YS(N659));
   FAX1 add_291_U1_14 ( .A(digest[142]),  .B(d_reg[14]),  .C(add_291_carry[14]), .YC(add_291_carry[15]), .YS(N660));
   FAX1 add_291_U1_15 ( .A(digest[143]),  .B(d_reg[15]),  .C(add_291_carry[15]), .YC(add_291_carry[16]), .YS(N661));
   FAX1 add_291_U1_16 ( .A(digest[144]),  .B(d_reg[16]),  .C(add_291_carry[16]), .YC(add_291_carry[17]), .YS(N662));
   FAX1 add_291_U1_17 ( .A(digest[145]),  .B(d_reg[17]),  .C(add_291_carry[17]), .YC(add_291_carry[18]), .YS(N663));
   FAX1 add_291_U1_18 ( .A(digest[146]),  .B(d_reg[18]),  .C(add_291_carry[18]), .YC(add_291_carry[19]), .YS(N664));
   FAX1 add_291_U1_19 ( .A(digest[147]),  .B(d_reg[19]),  .C(add_291_carry[19]), .YC(add_291_carry[20]), .YS(N665));
   FAX1 add_291_U1_20 ( .A(digest[148]),  .B(d_reg[20]),  .C(add_291_carry[20]), .YC(add_291_carry[21]), .YS(N666));
   FAX1 add_291_U1_21 ( .A(digest[149]),  .B(d_reg[21]),  .C(add_291_carry[21]), .YC(add_291_carry[22]), .YS(N667));
   FAX1 add_291_U1_22 ( .A(digest[150]),  .B(d_reg[22]),  .C(add_291_carry[22]), .YC(add_291_carry[23]), .YS(N668));
   FAX1 add_291_U1_23 ( .A(digest[151]),  .B(d_reg[23]),  .C(add_291_carry[23]), .YC(add_291_carry[24]), .YS(N669));
   FAX1 add_291_U1_24 ( .A(digest[152]),  .B(d_reg[24]),  .C(add_291_carry[24]), .YC(add_291_carry[25]), .YS(N670));
   FAX1 add_291_U1_25 ( .A(digest[153]),  .B(d_reg[25]),  .C(add_291_carry[25]), .YC(add_291_carry[26]), .YS(N671));
   FAX1 add_291_U1_26 ( .A(digest[154]),  .B(d_reg[26]),  .C(add_291_carry[26]), .YC(add_291_carry[27]), .YS(N672));
   FAX1 add_291_U1_27 ( .A(digest[155]),  .B(d_reg[27]),  .C(add_291_carry[27]), .YC(add_291_carry[28]), .YS(N673));
   FAX1 add_291_U1_28 ( .A(digest[156]),  .B(d_reg[28]),  .C(add_291_carry[28]), .YC(add_291_carry[29]), .YS(N674));
   FAX1 add_291_U1_29 ( .A(digest[157]),  .B(d_reg[29]),  .C(add_291_carry[29]), .YC(add_291_carry[30]), .YS(N675));
   FAX1 add_291_U1_30 ( .A(digest[158]),  .B(d_reg[30]),  .C(add_291_carry[30]), .YC(add_291_carry[31]), .YS(N676));
   FAX1 add_291_U1_31 ( .A(digest[159]),  .B(d_reg[31]),  .C(add_291_carry[31]), .YS(N677));
   FAX1 add_290_U1_1 ( .A(digest[161]),  .B(c_reg[1]),  .C(n2972), .YC(add_290_carry[2]), .YS(N615));
   FAX1 add_290_U1_2 ( .A(digest[162]),  .B(c_reg[2]),  .C(add_290_carry[2]), .YC(add_290_carry[3]), .YS(N616));
   FAX1 add_290_U1_3 ( .A(digest[163]),  .B(c_reg[3]),  .C(add_290_carry[3]), .YC(add_290_carry[4]), .YS(N617));
   FAX1 add_290_U1_4 ( .A(digest[164]),  .B(c_reg[4]),  .C(add_290_carry[4]), .YC(add_290_carry[5]), .YS(N618));
   FAX1 add_290_U1_5 ( .A(digest[165]),  .B(c_reg[5]),  .C(add_290_carry[5]), .YC(add_290_carry[6]), .YS(N619));
   FAX1 add_290_U1_6 ( .A(digest[166]),  .B(c_reg[6]),  .C(add_290_carry[6]), .YC(add_290_carry[7]), .YS(N620));
   FAX1 add_290_U1_7 ( .A(digest[167]),  .B(c_reg[7]),  .C(add_290_carry[7]), .YC(add_290_carry[8]), .YS(N621));
   FAX1 add_290_U1_8 ( .A(digest[168]),  .B(c_reg[8]),  .C(add_290_carry[8]), .YC(add_290_carry[9]), .YS(N622));
   FAX1 add_290_U1_9 ( .A(digest[169]),  .B(c_reg[9]),  .C(add_290_carry[9]), .YC(add_290_carry[10]), .YS(N623));
   FAX1 add_290_U1_10 ( .A(digest[170]),  .B(c_reg[10]),  .C(add_290_carry[10]), .YC(add_290_carry[11]), .YS(N624));
   FAX1 add_290_U1_11 ( .A(digest[171]),  .B(c_reg[11]),  .C(add_290_carry[11]), .YC(add_290_carry[12]), .YS(N625));
   FAX1 add_290_U1_12 ( .A(digest[172]),  .B(c_reg[12]),  .C(add_290_carry[12]), .YC(add_290_carry[13]), .YS(N626));
   FAX1 add_290_U1_13 ( .A(digest[173]),  .B(c_reg[13]),  .C(add_290_carry[13]), .YC(add_290_carry[14]), .YS(N627));
   FAX1 add_290_U1_14 ( .A(digest[174]),  .B(c_reg[14]),  .C(add_290_carry[14]), .YC(add_290_carry[15]), .YS(N628));
   FAX1 add_290_U1_15 ( .A(digest[175]),  .B(c_reg[15]),  .C(add_290_carry[15]), .YC(add_290_carry[16]), .YS(N629));
   FAX1 add_290_U1_16 ( .A(digest[176]),  .B(c_reg[16]),  .C(add_290_carry[16]), .YC(add_290_carry[17]), .YS(N630));
   FAX1 add_290_U1_17 ( .A(digest[177]),  .B(c_reg[17]),  .C(add_290_carry[17]), .YC(add_290_carry[18]), .YS(N631));
   FAX1 add_290_U1_18 ( .A(digest[178]),  .B(c_reg[18]),  .C(add_290_carry[18]), .YC(add_290_carry[19]), .YS(N632));
   FAX1 add_290_U1_19 ( .A(digest[179]),  .B(c_reg[19]),  .C(add_290_carry[19]), .YC(add_290_carry[20]), .YS(N633));
   FAX1 add_290_U1_20 ( .A(digest[180]),  .B(c_reg[20]),  .C(add_290_carry[20]), .YC(add_290_carry[21]), .YS(N634));
   FAX1 add_290_U1_21 ( .A(digest[181]),  .B(c_reg[21]),  .C(add_290_carry[21]), .YC(add_290_carry[22]), .YS(N635));
   FAX1 add_290_U1_22 ( .A(digest[182]),  .B(c_reg[22]),  .C(add_290_carry[22]), .YC(add_290_carry[23]), .YS(N636));
   FAX1 add_290_U1_23 ( .A(digest[183]),  .B(c_reg[23]),  .C(add_290_carry[23]), .YC(add_290_carry[24]), .YS(N637));
   FAX1 add_290_U1_24 ( .A(digest[184]),  .B(c_reg[24]),  .C(add_290_carry[24]), .YC(add_290_carry[25]), .YS(N638));
   FAX1 add_290_U1_25 ( .A(digest[185]),  .B(c_reg[25]),  .C(add_290_carry[25]), .YC(add_290_carry[26]), .YS(N639));
   FAX1 add_290_U1_26 ( .A(digest[186]),  .B(c_reg[26]),  .C(add_290_carry[26]), .YC(add_290_carry[27]), .YS(N640));
   FAX1 add_290_U1_27 ( .A(digest[187]),  .B(c_reg[27]),  .C(add_290_carry[27]), .YC(add_290_carry[28]), .YS(N641));
   FAX1 add_290_U1_28 ( .A(digest[188]),  .B(c_reg[28]),  .C(add_290_carry[28]), .YC(add_290_carry[29]), .YS(N642));
   FAX1 add_290_U1_29 ( .A(digest[189]),  .B(c_reg[29]),  .C(add_290_carry[29]), .YC(add_290_carry[30]), .YS(N643));
   FAX1 add_290_U1_30 ( .A(digest[190]),  .B(c_reg[30]),  .C(add_290_carry[30]), .YC(add_290_carry[31]), .YS(N644));
   FAX1 add_290_U1_31 ( .A(digest[191]),  .B(c_reg[31]),  .C(add_290_carry[31]), .YS(N645));
   FAX1 add_289_U1_1 ( .A(digest[193]),  .B(b_reg[1]),  .C(n2968), .YC(add_289_carry[2]), .YS(N583));
   FAX1 add_289_U1_2 ( .A(digest[194]),  .B(b_reg[2]),  .C(add_289_carry[2]), .YC(add_289_carry[3]), .YS(N584));
   FAX1 add_289_U1_3 ( .A(digest[195]),  .B(b_reg[3]),  .C(add_289_carry[3]), .YC(add_289_carry[4]), .YS(N585));
   FAX1 add_289_U1_4 ( .A(digest[196]),  .B(b_reg[4]),  .C(add_289_carry[4]), .YC(add_289_carry[5]), .YS(N586));
   FAX1 add_289_U1_5 ( .A(digest[197]),  .B(b_reg[5]),  .C(add_289_carry[5]), .YC(add_289_carry[6]), .YS(N587));
   FAX1 add_289_U1_6 ( .A(digest[198]),  .B(b_reg[6]),  .C(add_289_carry[6]), .YC(add_289_carry[7]), .YS(N588));
   FAX1 add_289_U1_7 ( .A(digest[199]),  .B(b_reg[7]),  .C(add_289_carry[7]), .YC(add_289_carry[8]), .YS(N589));
   FAX1 add_289_U1_8 ( .A(digest[200]),  .B(b_reg[8]),  .C(add_289_carry[8]), .YC(add_289_carry[9]), .YS(N590));
   FAX1 add_289_U1_9 ( .A(digest[201]),  .B(b_reg[9]),  .C(add_289_carry[9]), .YC(add_289_carry[10]), .YS(N591));
   FAX1 add_289_U1_10 ( .A(digest[202]),  .B(b_reg[10]),  .C(add_289_carry[10]), .YC(add_289_carry[11]), .YS(N592));
   FAX1 add_289_U1_11 ( .A(digest[203]),  .B(b_reg[11]),  .C(add_289_carry[11]), .YC(add_289_carry[12]), .YS(N593));
   FAX1 add_289_U1_12 ( .A(digest[204]),  .B(b_reg[12]),  .C(add_289_carry[12]), .YC(add_289_carry[13]), .YS(N594));
   FAX1 add_289_U1_13 ( .A(digest[205]),  .B(b_reg[13]),  .C(add_289_carry[13]), .YC(add_289_carry[14]), .YS(N595));
   FAX1 add_289_U1_14 ( .A(digest[206]),  .B(b_reg[14]),  .C(add_289_carry[14]), .YC(add_289_carry[15]), .YS(N596));
   FAX1 add_289_U1_15 ( .A(digest[207]),  .B(b_reg[15]),  .C(add_289_carry[15]), .YC(add_289_carry[16]), .YS(N597));
   FAX1 add_289_U1_16 ( .A(digest[208]),  .B(b_reg[16]),  .C(add_289_carry[16]), .YC(add_289_carry[17]), .YS(N598));
   FAX1 add_289_U1_17 ( .A(digest[209]),  .B(b_reg[17]),  .C(add_289_carry[17]), .YC(add_289_carry[18]), .YS(N599));
   FAX1 add_289_U1_18 ( .A(digest[210]),  .B(b_reg[18]),  .C(add_289_carry[18]), .YC(add_289_carry[19]), .YS(N600));
   FAX1 add_289_U1_19 ( .A(digest[211]),  .B(b_reg[19]),  .C(add_289_carry[19]), .YC(add_289_carry[20]), .YS(N601));
   FAX1 add_289_U1_20 ( .A(digest[212]),  .B(b_reg[20]),  .C(add_289_carry[20]), .YC(add_289_carry[21]), .YS(N602));
   FAX1 add_289_U1_21 ( .A(digest[213]),  .B(b_reg[21]),  .C(add_289_carry[21]), .YC(add_289_carry[22]), .YS(N603));
   FAX1 add_289_U1_22 ( .A(digest[214]),  .B(b_reg[22]),  .C(add_289_carry[22]), .YC(add_289_carry[23]), .YS(N604));
   FAX1 add_289_U1_23 ( .A(digest[215]),  .B(b_reg[23]),  .C(add_289_carry[23]), .YC(add_289_carry[24]), .YS(N605));
   FAX1 add_289_U1_24 ( .A(digest[216]),  .B(b_reg[24]),  .C(add_289_carry[24]), .YC(add_289_carry[25]), .YS(N606));
   FAX1 add_289_U1_25 ( .A(digest[217]),  .B(b_reg[25]),  .C(add_289_carry[25]), .YC(add_289_carry[26]), .YS(N607));
   FAX1 add_289_U1_26 ( .A(digest[218]),  .B(b_reg[26]),  .C(add_289_carry[26]), .YC(add_289_carry[27]), .YS(N608));
   FAX1 add_289_U1_27 ( .A(digest[219]),  .B(b_reg[27]),  .C(add_289_carry[27]), .YC(add_289_carry[28]), .YS(N609));
   FAX1 add_289_U1_28 ( .A(digest[220]),  .B(b_reg[28]),  .C(add_289_carry[28]), .YC(add_289_carry[29]), .YS(N610));
   FAX1 add_289_U1_29 ( .A(digest[221]),  .B(b_reg[29]),  .C(add_289_carry[29]), .YC(add_289_carry[30]), .YS(N611));
   FAX1 add_289_U1_30 ( .A(digest[222]),  .B(b_reg[30]),  .C(add_289_carry[30]), .YC(add_289_carry[31]), .YS(N612));
   FAX1 add_289_U1_31 ( .A(digest[223]),  .B(b_reg[31]),  .C(add_289_carry[31]), .YS(N613));
   FAX1 add_288_U1_1 ( .A(digest[225]),  .B(a_reg[1]),  .C(n2973), .YC(add_288_carry[2]), .YS(N551));
   FAX1 add_288_U1_2 ( .A(digest[226]),  .B(a_reg[2]),  .C(add_288_carry[2]), .YC(add_288_carry[3]), .YS(N552));
   FAX1 add_288_U1_3 ( .A(digest[227]),  .B(a_reg[3]),  .C(add_288_carry[3]), .YC(add_288_carry[4]), .YS(N553));
   FAX1 add_288_U1_4 ( .A(digest[228]),  .B(a_reg[4]),  .C(add_288_carry[4]), .YC(add_288_carry[5]), .YS(N554));
   FAX1 add_288_U1_5 ( .A(digest[229]),  .B(a_reg[5]),  .C(add_288_carry[5]), .YC(add_288_carry[6]), .YS(N555));
   FAX1 add_288_U1_6 ( .A(digest[230]),  .B(a_reg[6]),  .C(add_288_carry[6]), .YC(add_288_carry[7]), .YS(N556));
   FAX1 add_288_U1_7 ( .A(digest[231]),  .B(a_reg[7]),  .C(add_288_carry[7]), .YC(add_288_carry[8]), .YS(N557));
   FAX1 add_288_U1_8 ( .A(digest[232]),  .B(a_reg[8]),  .C(add_288_carry[8]), .YC(add_288_carry[9]), .YS(N558));
   FAX1 add_288_U1_9 ( .A(digest[233]),  .B(a_reg[9]),  .C(add_288_carry[9]), .YC(add_288_carry[10]), .YS(N559));
   FAX1 add_288_U1_10 ( .A(digest[234]),  .B(a_reg[10]),  .C(add_288_carry[10]), .YC(add_288_carry[11]), .YS(N560));
   FAX1 add_288_U1_11 ( .A(digest[235]),  .B(a_reg[11]),  .C(add_288_carry[11]), .YC(add_288_carry[12]), .YS(N561));
   FAX1 add_288_U1_12 ( .A(digest[236]),  .B(a_reg[12]),  .C(add_288_carry[12]), .YC(add_288_carry[13]), .YS(N562));
   FAX1 add_288_U1_13 ( .A(digest[237]),  .B(a_reg[13]),  .C(add_288_carry[13]), .YC(add_288_carry[14]), .YS(N563));
   FAX1 add_288_U1_14 ( .A(digest[238]),  .B(a_reg[14]),  .C(add_288_carry[14]), .YC(add_288_carry[15]), .YS(N564));
   FAX1 add_288_U1_15 ( .A(digest[239]),  .B(a_reg[15]),  .C(add_288_carry[15]), .YC(add_288_carry[16]), .YS(N565));
   FAX1 add_288_U1_16 ( .A(digest[240]),  .B(a_reg[16]),  .C(add_288_carry[16]), .YC(add_288_carry[17]), .YS(N566));
   FAX1 add_288_U1_17 ( .A(digest[241]),  .B(a_reg[17]),  .C(add_288_carry[17]), .YC(add_288_carry[18]), .YS(N567));
   FAX1 add_288_U1_18 ( .A(digest[242]),  .B(a_reg[18]),  .C(add_288_carry[18]), .YC(add_288_carry[19]), .YS(N568));
   FAX1 add_288_U1_19 ( .A(digest[243]),  .B(a_reg[19]),  .C(add_288_carry[19]), .YC(add_288_carry[20]), .YS(N569));
   FAX1 add_288_U1_20 ( .A(digest[244]),  .B(a_reg[20]),  .C(add_288_carry[20]), .YC(add_288_carry[21]), .YS(N570));
   FAX1 add_288_U1_21 ( .A(digest[245]),  .B(a_reg[21]),  .C(add_288_carry[21]), .YC(add_288_carry[22]), .YS(N571));
   FAX1 add_288_U1_22 ( .A(digest[246]),  .B(a_reg[22]),  .C(add_288_carry[22]), .YC(add_288_carry[23]), .YS(N572));
   FAX1 add_288_U1_23 ( .A(digest[247]),  .B(a_reg[23]),  .C(add_288_carry[23]), .YC(add_288_carry[24]), .YS(N573));
   FAX1 add_288_U1_24 ( .A(digest[248]),  .B(a_reg[24]),  .C(add_288_carry[24]), .YC(add_288_carry[25]), .YS(N574));
   FAX1 add_288_U1_25 ( .A(digest[249]),  .B(a_reg[25]),  .C(add_288_carry[25]), .YC(add_288_carry[26]), .YS(N575));
   FAX1 add_288_U1_26 ( .A(digest[250]),  .B(a_reg[26]),  .C(add_288_carry[26]), .YC(add_288_carry[27]), .YS(N576));
   FAX1 add_288_U1_27 ( .A(digest[251]),  .B(a_reg[27]),  .C(add_288_carry[27]), .YC(add_288_carry[28]), .YS(N577));
   FAX1 add_288_U1_28 ( .A(digest[252]),  .B(a_reg[28]),  .C(add_288_carry[28]), .YC(add_288_carry[29]), .YS(N578));
   FAX1 add_288_U1_29 ( .A(digest[253]),  .B(a_reg[29]),  .C(add_288_carry[29]), .YC(add_288_carry[30]), .YS(N579));
   FAX1 add_288_U1_30 ( .A(digest[254]),  .B(a_reg[30]),  .C(add_288_carry[30]), .YC(add_288_carry[31]), .YS(N580));
   FAX1 add_288_U1_31 ( .A(digest[255]),  .B(a_reg[31]),  .C(add_288_carry[31]), .YS(N581));
   AND2X1 U1851 ( .A(n2718),  .B(n2595), .Y(n5971));
   AND2X1 U1852 ( .A(n5821),  .B(n2893), .Y(n5991));
   AND2X1 U1853 ( .A(n2847),  .B(n2783), .Y(n5770));
   AND2X1 U1854 ( .A(n2657),  .B(n2720), .Y(n5751));
   AND2X1 U1855 ( .A(n2890),  .B(n2107), .Y(n5749));
   AND2X1 U1856 ( .A(n2847),  .B(n2845), .Y(n6033));
   AND2X1 U1857 ( .A(n5839),  .B(n2712), .Y(n5837));
   AND2X1 U1858 ( .A(n2894),  .B(n2958), .Y(n4169));
   AND2X1 U1859 ( .A(n2955),  .B(n2717), .Y(n5853));
   AND2X1 U1860 ( .A(n4442),  .B(n1953), .Y(n4170));
   AND2X1 U1861 ( .A(n5771),  .B(n2955), .Y(n5752));
   AND2X1 U1862 ( .A(n5786),  .B(n2720), .Y(n5793));
   OR2X1 U1863 ( .A(n2717),  .B(n5843), .Y(n5867));
   AND2X1 U1864 ( .A(n2777),  .B(n3100), .Y(n3103));
   OR2X1 U1865 ( .A(n5912),  .B(n1777), .Y(n1756));
   OR2X1 U1866 ( .A(n2023),  .B(n1778), .Y(n1757));
   OR2X1 U1867 ( .A(n2100),  .B(n1776), .Y(n1758));
   AND2X1 U1868 ( .A(n2951),  .B(n4713), .Y(n4783));
   OR2X1 U1869 ( .A(n2127),  .B(n1780), .Y(n1759));
   OR2X1 U1870 ( .A(n2065),  .B(n1866), .Y(n1760));
   OR2X1 U1871 ( .A(n2068),  .B(n1867), .Y(n1761));
   OR2X1 U1872 ( .A(n2071),  .B(n1858), .Y(n1762));
   OR2X1 U1873 ( .A(n2074),  .B(n1856), .Y(n1763));
   OR2X1 U1874 ( .A(n2077),  .B(n1859), .Y(n1764));
   OR2X1 U1875 ( .A(n2082),  .B(n1860), .Y(n1765));
   OR2X1 U1876 ( .A(n2085),  .B(n1865), .Y(n1766));
   OR2X1 U1877 ( .A(n2091),  .B(n1868), .Y(n1767));
   OR2X1 U1878 ( .A(n2094),  .B(n1869), .Y(n1768));
   OR2X1 U1879 ( .A(n2046),  .B(n1861), .Y(n1769));
   OR2X1 U1880 ( .A(n2048),  .B(n1855), .Y(n1770));
   OR2X1 U1881 ( .A(n2051),  .B(n1862), .Y(n1771));
   OR2X1 U1882 ( .A(n2054),  .B(n1863), .Y(n1772));
   OR2X1 U1883 ( .A(n2057),  .B(n1864), .Y(n1773));
   OR2X1 U1884 ( .A(n2062),  .B(n1857), .Y(n1774));
   AND2X1 U1885 ( .A(n2891),  .B(n2720), .Y(n5848));
   AND2X1 U1886 ( .A(n2849),  .B(n2720), .Y(n5861));
   OR2X1 U1887 ( .A(n1936),  .B(n1854), .Y(n1775));
   OR2X1 U1888 ( .A(n2099),  .B(n1871), .Y(n1776));
   OR2X1 U1889 ( .A(n1877),  .B(n5981), .Y(n1777));
   OR2X1 U1890 ( .A(n1898),  .B(n2022), .Y(n1778));
   OR2X1 U1891 ( .A(n1941),  .B(n1875), .Y(n1779));
   OR2X1 U1892 ( .A(n3115),  .B(rst), .Y(n1780));
   OR2X1 U1893 ( .A(n1974),  .B(n1872), .Y(n1781));
   OR2X1 U1894 ( .A(n1878),  .B(n1982), .Y(n1782));
   OR2X1 U1895 ( .A(n1879),  .B(n1984), .Y(n1783));
   OR2X1 U1896 ( .A(n1880),  .B(n1986), .Y(n1784));
   OR2X1 U1897 ( .A(n1881),  .B(n1988), .Y(n1785));
   OR2X1 U1898 ( .A(n1882),  .B(n1990), .Y(n1786));
   OR2X1 U1899 ( .A(n1883),  .B(n1992), .Y(n1787));
   OR2X1 U1900 ( .A(n1884),  .B(n1994), .Y(n1788));
   OR2X1 U1901 ( .A(n1885),  .B(n1996), .Y(n1789));
   OR2X1 U1902 ( .A(n1886),  .B(n1998), .Y(n1790));
   OR2X1 U1903 ( .A(n1887),  .B(n2000), .Y(n1791));
   OR2X1 U1904 ( .A(n1888),  .B(n2002), .Y(n1792));
   OR2X1 U1905 ( .A(n1889),  .B(n2004), .Y(n1793));
   OR2X1 U1906 ( .A(n1890),  .B(n2006), .Y(n1794));
   OR2X1 U1907 ( .A(n1891),  .B(n2008), .Y(n1795));
   OR2X1 U1908 ( .A(n1892),  .B(n2010), .Y(n1796));
   OR2X1 U1909 ( .A(n1893),  .B(n2012), .Y(n1797));
   OR2X1 U1910 ( .A(n1894),  .B(n2014), .Y(n1798));
   OR2X1 U1911 ( .A(n1895),  .B(n2016), .Y(n1799));
   OR2X1 U1912 ( .A(n1896),  .B(n2018), .Y(n1800));
   OR2X1 U1913 ( .A(n1897),  .B(n2020), .Y(n1801));
   OR2X1 U1914 ( .A(n1899),  .B(n2024), .Y(n1802));
   OR2X1 U1915 ( .A(n1900),  .B(n2026), .Y(n1803));
   OR2X1 U1916 ( .A(n1901),  .B(n2028), .Y(n1804));
   OR2X1 U1917 ( .A(n1902),  .B(n2030), .Y(n1805));
   OR2X1 U1918 ( .A(n1903),  .B(n2032), .Y(n1806));
   OR2X1 U1919 ( .A(n1904),  .B(n2034), .Y(n1807));
   OR2X1 U1920 ( .A(n1905),  .B(n2036), .Y(n1808));
   OR2X1 U1921 ( .A(n1906),  .B(n2038), .Y(n1809));
   OR2X1 U1922 ( .A(n1907),  .B(n2040), .Y(n1810));
   OR2X1 U1923 ( .A(n1908),  .B(n2042), .Y(n1811));
   OR2X1 U1924 ( .A(n1876),  .B(n2095), .Y(n1812));
   OR2X1 U1925 ( .A(n1874),  .B(n2078), .Y(n1813));
   OR2X1 U1926 ( .A(n1873),  .B(n2087), .Y(n1814));
   OR2X1 U1927 ( .A(n2058),  .B(n1870), .Y(n1815));
   OR2X1 U1928 ( .A(n2059),  .B(n1815), .Y(n1816));
   OR2X1 U1929 ( .A(n2088),  .B(n1814), .Y(n1817));
   OR2X1 U1930 ( .A(n2079),  .B(n1813), .Y(n1818));
   OR2X1 U1931 ( .A(n2019),  .B(n1800), .Y(n1819));
   OR2X1 U1932 ( .A(n2021),  .B(n1801), .Y(n1820));
   OR2X1 U1933 ( .A(n2025),  .B(n1802), .Y(n1821));
   OR2X1 U1934 ( .A(n2027),  .B(n1803), .Y(n1822));
   OR2X1 U1935 ( .A(n2029),  .B(n1804), .Y(n1823));
   OR2X1 U1936 ( .A(n2031),  .B(n1805), .Y(n1824));
   OR2X1 U1937 ( .A(n2033),  .B(n1806), .Y(n1825));
   OR2X1 U1938 ( .A(n2035),  .B(n1807), .Y(n1826));
   OR2X1 U1939 ( .A(n2037),  .B(n1808), .Y(n1827));
   OR2X1 U1940 ( .A(n2039),  .B(n1809), .Y(n1828));
   OR2X1 U1941 ( .A(n2041),  .B(n1810), .Y(n1829));
   OR2X1 U1942 ( .A(n2043),  .B(n1811), .Y(n1830));
   OR2X1 U1943 ( .A(n1997),  .B(n1789), .Y(n1831));
   OR2X1 U1944 ( .A(n1999),  .B(n1790), .Y(n1832));
   OR2X1 U1945 ( .A(n2003),  .B(n1792), .Y(n1833));
   OR2X1 U1946 ( .A(n2005),  .B(n1793), .Y(n1834));
   OR2X1 U1947 ( .A(n2007),  .B(n1794), .Y(n1835));
   OR2X1 U1948 ( .A(n2009),  .B(n1795), .Y(n1836));
   OR2X1 U1949 ( .A(n2011),  .B(n1796), .Y(n1837));
   OR2X1 U1950 ( .A(n2013),  .B(n1797), .Y(n1838));
   OR2X1 U1951 ( .A(n2015),  .B(n1798), .Y(n1839));
   OR2X1 U1952 ( .A(n2017),  .B(n1799), .Y(n1840));
   OR2X1 U1953 ( .A(n1983),  .B(n1782), .Y(n1841));
   OR2X1 U1954 ( .A(n1985),  .B(n1783), .Y(n1842));
   OR2X1 U1955 ( .A(n1987),  .B(n1784), .Y(n1843));
   OR2X1 U1956 ( .A(n1989),  .B(n1785), .Y(n1844));
   OR2X1 U1957 ( .A(n1991),  .B(n1786), .Y(n1845));
   OR2X1 U1958 ( .A(n1993),  .B(n1787), .Y(n1846));
   OR2X1 U1959 ( .A(n1995),  .B(n1788), .Y(n1847));
   OR2X1 U1960 ( .A(n2001),  .B(n1791), .Y(n1848));
   OR2X1 U1961 ( .A(n2096),  .B(n1812), .Y(n1849));
   AND2X1 U1962 ( .A(n1849),  .B(N869), .Y(n1850));
   OR2X1 U1963 ( .A(n1975),  .B(n1781), .Y(n1851));
   AND2X1 U1964 ( .A(n2891),  .B(n2657), .Y(n5786));
   AND2X1 U1965 ( .A(n2849),  .B(n2657), .Y(n5816));
   OR2X1 U1966 ( .A(n3116),  .B(rst), .Y(n1852));
   OR2X1 U1967 ( .A(n1942),  .B(n1779), .Y(n1853));
   AND2X1 U1968 ( .A(n2782),  .B(n2098), .Y(n5849));
   OR2X1 U1969 ( .A(n1935),  .B(n1756), .Y(n1854));
   OR2X1 U1970 ( .A(n2047),  .B(n1758), .Y(n1855));
   OR2X1 U1971 ( .A(n2073),  .B(n1969), .Y(n1856));
   OR2X1 U1972 ( .A(n2060),  .B(n2061), .Y(n1857));
   OR2X1 U1973 ( .A(n2069),  .B(n2070), .Y(n1858));
   OR2X1 U1974 ( .A(n2075),  .B(n2076), .Y(n1859));
   OR2X1 U1975 ( .A(n2080),  .B(n2081), .Y(n1860));
   OR2X1 U1976 ( .A(n2044),  .B(n2045), .Y(n1861));
   OR2X1 U1977 ( .A(n2049),  .B(n2050), .Y(n1862));
   OR2X1 U1978 ( .A(n2052),  .B(n2053), .Y(n1863));
   OR2X1 U1979 ( .A(n2055),  .B(n2056), .Y(n1864));
   OR2X1 U1980 ( .A(n2083),  .B(n2084), .Y(n1865));
   OR2X1 U1981 ( .A(n2063),  .B(n2064), .Y(n1866));
   OR2X1 U1982 ( .A(n2066),  .B(n2067), .Y(puf_1_wire_3));
   OR2X1 U1983 ( .A(n2089),  .B(n2090), .Y(n1868));
   OR2X1 U1984 ( .A(n2092),  .B(n2093), .Y(n1869));
   AND2X1 U1985 ( .A(n5845),  .B(n5917), .Y(n1870));
   AND2X1 U1986 ( .A(n5782),  .B(n2785), .Y(n1871));
   AND2X1 U1987 ( .A(n5771),  .B(n2719), .Y(n1872));
   OR2X2 U1988 ( .A(n6064),  .B(n6065), .Y(n1873));
   OR2X2 U1989 ( .A(n5996),  .B(n5997), .Y(n1874));
   AND2X1 U1990 ( .A(n5886),  .B(n2591), .Y(n1875));
   AND2X1 U1991 ( .A(w_mem_inst_w_new[0]),  .B(n2957), .Y(n1876));
   AND2X1 U1992 ( .A(n5936),  .B(n5789), .Y(n1877));
   AND2X1 U1993 ( .A(w_mem_inst_w_new[9]),  .B(n2957), .Y(n1878));
   AND2X1 U1994 ( .A(w_mem_inst_w_new[8]),  .B(n2957), .Y(n1879));
   AND2X1 U1995 ( .A(w_mem_inst_w_new[7]),  .B(n2957), .Y(n1880));
   AND2X1 U1996 ( .A(w_mem_inst_w_new[6]),  .B(n2957), .Y(n1881));
   AND2X1 U1997 ( .A(w_mem_inst_w_new[5]),  .B(n2957), .Y(n1882));
   AND2X1 U1998 ( .A(w_mem_inst_w_new[4]),  .B(n2957), .Y(n1883));
   AND2X1 U1999 ( .A(w_mem_inst_w_new[3]),  .B(n2957), .Y(n1884));
   AND2X1 U2000 ( .A(w_mem_inst_w_new[31]),  .B(n2957), .Y(n1885));
   AND2X1 U2001 ( .A(w_mem_inst_w_new[30]),  .B(n2957), .Y(n1886));
   AND2X1 U2002 ( .A(w_mem_inst_w_new[2]),  .B(n2957), .Y(n1887));
   AND2X1 U2003 ( .A(w_mem_inst_w_new[29]),  .B(n2957), .Y(n1888));
   AND2X1 U2004 ( .A(w_mem_inst_w_new[28]),  .B(n2957), .Y(n1889));
   AND2X1 U2005 ( .A(w_mem_inst_w_new[27]),  .B(n2957), .Y(n1890));
   AND2X1 U2006 ( .A(w_mem_inst_w_new[26]),  .B(n2957), .Y(n1891));
   AND2X1 U2007 ( .A(w_mem_inst_w_new[25]),  .B(n2957), .Y(n1892));
   AND2X1 U2008 ( .A(w_mem_inst_w_new[24]),  .B(n2957), .Y(n1893));
   AND2X1 U2009 ( .A(w_mem_inst_w_new[23]),  .B(n2957), .Y(n1894));
   AND2X1 U2010 ( .A(w_mem_inst_w_new[22]),  .B(n2957), .Y(n1895));
   AND2X1 U2011 ( .A(w_mem_inst_w_new[21]),  .B(n2957), .Y(n1896));
   AND2X1 U2012 ( .A(w_mem_inst_w_new[20]),  .B(n2957), .Y(n1897));
   AND2X1 U2013 ( .A(w_mem_inst_w_new[1]),  .B(n2957), .Y(n1898));
   AND2X1 U2014 ( .A(w_mem_inst_w_new[19]),  .B(n2957), .Y(n1899));
   AND2X1 U2015 ( .A(w_mem_inst_w_new[18]),  .B(n2957), .Y(n1900));
   AND2X1 U2016 ( .A(w_mem_inst_w_new[17]),  .B(n2957), .Y(n1901));
   AND2X1 U2017 ( .A(w_mem_inst_w_new[16]),  .B(n2957), .Y(n1902));
   AND2X1 U2018 ( .A(w_mem_inst_w_new[15]),  .B(n2957), .Y(n1903));
   AND2X1 U2019 ( .A(w_mem_inst_w_new[14]),  .B(n2957), .Y(n1904));
   AND2X1 U2020 ( .A(w_mem_inst_w_new[13]),  .B(n2957), .Y(n1905));
   AND2X1 U2021 ( .A(w_mem_inst_w_new[12]),  .B(n2957), .Y(n1906));
   AND2X1 U2022 ( .A(w_mem_inst_w_new[11]),  .B(n2957), .Y(n1907));
   AND2X1 U2023 ( .A(w_mem_inst_w_new[10]),  .B(n2957), .Y(n1908));
   BUFX2 U2024 ( .A(n5643), .Y(n1909));
   BUFX2 U2025 ( .A(n5647), .Y(n1910));
   BUFX2 U2026 ( .A(n5649), .Y(n1911));
   BUFX2 U2027 ( .A(n5651), .Y(n1912));
   BUFX2 U2028 ( .A(n5655), .Y(n1913));
   BUFX2 U2029 ( .A(n5657), .Y(n1914));
   BUFX2 U2030 ( .A(n5665), .Y(n1915));
   BUFX2 U2031 ( .A(n5667), .Y(n1916));
   BUFX2 U2032 ( .A(n5669), .Y(n1917));
   BUFX2 U2033 ( .A(n5671), .Y(n1918));
   BUFX2 U2034 ( .A(n5798), .Y(n1919));
   BUFX2 U2035 ( .A(n5804), .Y(n1920));
   BUFX2 U2036 ( .A(n5866), .Y(n1921));
   BUFX2 U2037 ( .A(n5871), .Y(n1922));
   BUFX2 U2038 ( .A(n5975), .Y(n1923));
   BUFX2 U2039 ( .A(n6012), .Y(n1924));
   BUFX2 U2040 ( .A(n6032), .Y(n1925));
   BUFX2 U2041 ( .A(n6035), .Y(n1926));
   BUFX2 U2042 ( .A(n6009), .Y(n1927));
   BUFX2 U2043 ( .A(n6081), .Y(n1928));
   BUFX2 U2044 ( .A(n6115), .Y(n1929));
   AND2X1 U2045 ( .A(t_ctr_reg[3]),  .B(n6000), .Y(n5780));
   INVX1 U2046 ( .A(n5780), .Y(n1930));
   AND2X1 U2047 ( .A(n5846),  .B(t_ctr_reg[4]), .Y(n5844));
   INVX1 U2048 ( .A(n5844), .Y(n1931));
   AND2X1 U2049 ( .A(n5874),  .B(n4707), .Y(n5890));
   INVX1 U2050 ( .A(n5890), .Y(n1932));
   AND2X1 U2051 ( .A(n6061),  .B(n4703), .Y(n6014));
   INVX1 U2052 ( .A(n6014), .Y(n1933));
   AND2X1 U2053 ( .A(n5814),  .B(n4705), .Y(n6039));
   INVX1 U2054 ( .A(n6039), .Y(n1934));
   INVX1 U2055 ( .A(n5785), .Y(n1935));
   INVX1 U2056 ( .A(n5784), .Y(n1936));
   BUFX2 U2057 ( .A(n5879), .Y(n1937));
   BUFX2 U2058 ( .A(n5946), .Y(n1938));
   BUFX2 U2059 ( .A(n6018), .Y(n1939));
   BUFX2 U2060 ( .A(n6059), .Y(n1940));
   INVX1 U2061 ( .A(n6091), .Y(n1941));
   INVX1 U2062 ( .A(n6090), .Y(n1942));
   BUFX2 U2063 ( .A(n6107), .Y(n1943));
   BUFX2 U2064 ( .A(n6122), .Y(n1944));
   BUFX2 U2065 ( .A(n5776), .Y(n1945));
   BUFX2 U2066 ( .A(n6019), .Y(n1946));
   BUFX2 U2067 ( .A(n6086), .Y(n1947));
   AND2X1 U2068 ( .A(n6061),  .B(n5763), .Y(n5981));
   BUFX2 U2069 ( .A(n5777), .Y(n1948));
   BUFX2 U2070 ( .A(n6020), .Y(n1949));
   BUFX2 U2071 ( .A(n6044), .Y(n1950));
   BUFX2 U2072 ( .A(n6087), .Y(n1951));
   BUFX2 U2073 ( .A(n6108), .Y(n1952));
   BUFX2 U2074 ( .A(n4663), .Y(n1953));
   BUFX2 U2075 ( .A(n5801), .Y(n1954));
   AND2X1 U2076 ( .A(n5814),  .B(n5789), .Y(n6067));
   INVX1 U2077 ( .A(n6067), .Y(n1955));
   BUFX2 U2078 ( .A(n6071), .Y(n1956));
   AND2X1 U2079 ( .A(n4703),  .B(n4707), .Y(n5788));
   INVX1 U2080 ( .A(n5788), .Y(n1957));
   AND2X1 U2081 ( .A(sha256_ctrl_reg[0]),  .B(n4692), .Y(n3115));
   INVX1 U2082 ( .A(n3115), .Y(n1958));
   AND2X1 U2083 ( .A(n2892),  .B(n2718), .Y(n5949));
   INVX1 U2084 ( .A(n5949), .Y(n1959));
   AND2X1 U2085 ( .A(n2782),  .B(n2953), .Y(n5915));
   INVX1 U2086 ( .A(n5915), .Y(n1960));
   BUFX2 U2087 ( .A(n5865), .Y(n1961));
   AND2X1 U2088 ( .A(n5763),  .B(n6000), .Y(n5803));
   INVX1 U2089 ( .A(n5803), .Y(n1962));
   AND2X1 U2090 ( .A(n2097),  .B(n2115), .Y(n5820));
   INVX1 U2091 ( .A(n5820), .Y(n1963));
   AND2X1 U2092 ( .A(n5917),  .B(n6000), .Y(n6050));
   INVX1 U2093 ( .A(n6050), .Y(n1964));
   BUFX2 U2094 ( .A(n5773), .Y(n1965));
   AND2X1 U2095 ( .A(n6000),  .B(n2785), .Y(n5783));
   INVX1 U2096 ( .A(n5783), .Y(n1966));
   AND2X1 U2097 ( .A(n5763),  .B(n6021), .Y(n6069));
   INVX1 U2098 ( .A(n6069), .Y(n1967));
   AND2X1 U2099 ( .A(n5846),  .B(n5789), .Y(n6003));
   INVX1 U2100 ( .A(n6003), .Y(n1968));
   BUFX2 U2101 ( .A(n5960), .Y(n1969));
   AND2X1 U2102 ( .A(n2890),  .B(n2714), .Y(n6024));
   INVX1 U2103 ( .A(n6024), .Y(n1970));
   AND2X1 U2104 ( .A(n6045),  .B(n4703), .Y(n6080));
   INVX1 U2105 ( .A(n6080), .Y(n1971));
   AND2X1 U2106 ( .A(n2954),  .B(n2097), .Y(n5799));
   INVX1 U2107 ( .A(n5799), .Y(n1972));
   AND2X1 U2108 ( .A(n2781),  .B(n2595), .Y(n5756));
   INVX1 U2109 ( .A(n5756), .Y(n1973));
   INVX1 U2110 ( .A(n6073), .Y(n1974));
   INVX1 U2111 ( .A(n6072), .Y(n1975));
   BUFX2 U2112 ( .A(n5812), .Y(n1976));
   AND2X1 U2113 ( .A(n2655),  .B(n2783), .Y(n5791));
   INVX1 U2114 ( .A(n5791), .Y(n1977));
   AND2X1 U2115 ( .A(n2718),  .B(n2651), .Y(n5750));
   INVX1 U2116 ( .A(n5750), .Y(n1978));
   AND2X1 U2117 ( .A(n2715),  .B(n2844), .Y(n5938));
   INVX1 U2118 ( .A(n5938), .Y(n1979));
   AND2X1 U2119 ( .A(n2116),  .B(n2115), .Y(n5830));
   INVX1 U2120 ( .A(n5830), .Y(n1980));
   AND2X1 U2121 ( .A(n2718),  .B(n2116), .Y(n5847));
   INVX1 U2122 ( .A(n5847), .Y(n1981));
   INVX1 U2123 ( .A(n4146), .Y(n1982));
   INVX1 U2124 ( .A(n4145), .Y(n1983));
   OR2X2 U2125 ( .A(n4147),  .B(n4148), .Y(n4146));
   INVX1 U2126 ( .A(n4173), .Y(n1984));
   INVX1 U2127 ( .A(n4172), .Y(n1985));
   OR2X2 U2128 ( .A(n4174),  .B(n4175), .Y(n4173));
   INVX1 U2129 ( .A(n4189), .Y(n1986));
   INVX1 U2130 ( .A(n4188), .Y(n1987));
   OR2X2 U2131 ( .A(n4190),  .B(n4191), .Y(n4189));
   INVX1 U2132 ( .A(n4205), .Y(n1988));
   INVX1 U2133 ( .A(n4204), .Y(n1989));
   OR2X2 U2134 ( .A(n4206),  .B(n4207), .Y(n4205));
   INVX1 U2135 ( .A(n4221), .Y(n1990));
   INVX1 U2136 ( .A(n4220), .Y(n1991));
   OR2X2 U2137 ( .A(n4222),  .B(n4223), .Y(n4221));
   INVX1 U2138 ( .A(n4237), .Y(n1992));
   INVX1 U2139 ( .A(n4236), .Y(n1993));
   OR2X2 U2140 ( .A(n4238),  .B(n4239), .Y(n4237));
   INVX1 U2141 ( .A(n4253), .Y(n1994));
   INVX1 U2142 ( .A(n4252), .Y(n1995));
   OR2X2 U2143 ( .A(n4254),  .B(n4255), .Y(n4253));
   INVX1 U2144 ( .A(n4269), .Y(n1996));
   INVX1 U2145 ( .A(n4268), .Y(n1997));
   OR2X2 U2146 ( .A(n4270),  .B(n4271), .Y(n4269));
   INVX1 U2147 ( .A(n4285), .Y(n1998));
   INVX1 U2148 ( .A(n4284), .Y(n1999));
   OR2X2 U2149 ( .A(n4286),  .B(n4287), .Y(n4285));
   INVX1 U2150 ( .A(n4301), .Y(n2000));
   INVX1 U2151 ( .A(n4300), .Y(n2001));
   OR2X2 U2152 ( .A(n4302),  .B(n4303), .Y(n4301));
   INVX1 U2153 ( .A(n4317), .Y(n2002));
   INVX1 U2154 ( .A(n4316), .Y(n2003));
   OR2X2 U2155 ( .A(n4318),  .B(n4319), .Y(n4317));
   INVX1 U2156 ( .A(n4333), .Y(n2004));
   INVX1 U2157 ( .A(n4332), .Y(n2005));
   OR2X2 U2158 ( .A(n4334),  .B(n4335), .Y(n4333));
   INVX1 U2159 ( .A(n4349), .Y(puf_2_wire_3));
   INVX1 U2160 ( .A(n4348), .Y(n2007));
   OR2X2 U2161 ( .A(n4350),  .B(n4351), .Y(n4349));
   INVX1 U2162 ( .A(n4365), .Y(n2008));
   INVX1 U2163 ( .A(n4364), .Y(n2009));
   OR2X2 U2164 ( .A(n4366),  .B(n4367), .Y(n4365));
   INVX1 U2165 ( .A(n4381), .Y(n2010));
   INVX1 U2166 ( .A(n4380), .Y(n2011));
   OR2X2 U2167 ( .A(n4382),  .B(n4383), .Y(n4381));
   INVX1 U2168 ( .A(n4397), .Y(n2012));
   INVX1 U2169 ( .A(n4396), .Y(n2013));
   OR2X2 U2170 ( .A(n4398),  .B(n4399), .Y(n4397));
   INVX1 U2171 ( .A(n4413), .Y(n2014));
   INVX1 U2172 ( .A(n4412), .Y(n2015));
   OR2X2 U2173 ( .A(n4414),  .B(n4415), .Y(n4413));
   INVX1 U2174 ( .A(n4429), .Y(n2016));
   INVX1 U2175 ( .A(n4428), .Y(n2017));
   OR2X2 U2176 ( .A(n4430),  .B(n4431), .Y(n4429));
   INVX1 U2177 ( .A(n4447), .Y(n2018));
   INVX1 U2178 ( .A(n4446), .Y(n2019));
   OR2X2 U2179 ( .A(n4448),  .B(n4449), .Y(n4447));
   INVX1 U2180 ( .A(n4463), .Y(n2020));
   INVX1 U2181 ( .A(n4462), .Y(n2021));
   OR2X2 U2182 ( .A(n4464),  .B(n4465), .Y(n4463));
   INVX1 U2183 ( .A(n4479), .Y(n2022));
   INVX1 U2184 ( .A(n4478), .Y(n2023));
   OR2X2 U2185 ( .A(n4480),  .B(n4481), .Y(n4479));
   INVX1 U2186 ( .A(n4495), .Y(n2024));
   INVX1 U2187 ( .A(n4494), .Y(n2025));
   OR2X2 U2188 ( .A(n4496),  .B(n4497), .Y(n4495));
   INVX1 U2189 ( .A(n4511), .Y(n2026));
   INVX1 U2190 ( .A(n4510), .Y(n2027));
   OR2X2 U2191 ( .A(n4512),  .B(n4513), .Y(n4511));
   INVX1 U2192 ( .A(n4527), .Y(n2028));
   INVX1 U2193 ( .A(n4526), .Y(n2029));
   OR2X2 U2194 ( .A(n4528),  .B(n4529), .Y(n4527));
   INVX1 U2195 ( .A(n4543), .Y(n2030));
   INVX1 U2196 ( .A(n4542), .Y(n2031));
   OR2X2 U2197 ( .A(n4544),  .B(n4545), .Y(n4543));
   INVX1 U2198 ( .A(n4559), .Y(n2032));
   INVX1 U2199 ( .A(n4558), .Y(n2033));
   OR2X2 U2200 ( .A(n4560),  .B(n4561), .Y(n4559));
   INVX1 U2201 ( .A(n4575), .Y(n2034));
   INVX1 U2202 ( .A(n4574), .Y(n2035));
   OR2X2 U2203 ( .A(n4576),  .B(n4577), .Y(n4575));
   INVX1 U2204 ( .A(n4591), .Y(n2036));
   INVX1 U2205 ( .A(n4590), .Y(n2037));
   OR2X2 U2206 ( .A(n4592),  .B(n4593), .Y(n4591));
   INVX1 U2207 ( .A(n4607), .Y(n2038));
   INVX1 U2208 ( .A(n4606), .Y(n2039));
   OR2X2 U2209 ( .A(n4608),  .B(n4609), .Y(n4607));
   INVX1 U2210 ( .A(n4623), .Y(n2040));
   INVX1 U2211 ( .A(n4622), .Y(n2041));
   OR2X2 U2212 ( .A(n4624),  .B(n4625), .Y(n4623));
   INVX1 U2213 ( .A(n4639), .Y(n2042));
   INVX1 U2214 ( .A(n4638), .Y(n2043));
   OR2X2 U2215 ( .A(n4640),  .B(n4641), .Y(n4639));
   INVX1 U2216 ( .A(n5744), .Y(n2044));
   INVX1 U2217 ( .A(n5743), .Y(n2045));
   INVX1 U2218 ( .A(n5742), .Y(n2046));
   INVX1 U2219 ( .A(n5759), .Y(n2047));
   INVX1 U2220 ( .A(n5758), .Y(n2048));
   INVX1 U2221 ( .A(n5810), .Y(n2049));
   INVX1 U2222 ( .A(n5809), .Y(n2050));
   INVX1 U2223 ( .A(n5808), .Y(n2051));
   INVX1 U2224 ( .A(n5825), .Y(n2052));
   INVX1 U2225 ( .A(n5824), .Y(n2053));
   INVX1 U2226 ( .A(n5823), .Y(n2054));
   INVX1 U2227 ( .A(n5835), .Y(n2055));
   INVX1 U2228 ( .A(n5834), .Y(n2056));
   INVX1 U2229 ( .A(n5833), .Y(n2057));
   INVX1 U2230 ( .A(n5851), .Y(n2058));
   INVX1 U2231 ( .A(n5850), .Y(n2059));
   INVX1 U2232 ( .A(n5878), .Y(n2060));
   INVX1 U2233 ( .A(n5877), .Y(n2061));
   INVX1 U2234 ( .A(n5876), .Y(n2062));
   INVX1 U2235 ( .A(n5907), .Y(n2063));
   INVX1 U2236 ( .A(n5906), .Y(n2064));
   INVX1 U2237 ( .A(n5905), .Y(n2065));
   AND2X2 U2238 ( .A(n5908),  .B(n5909), .Y(n5907));
   INVX1 U2239 ( .A(n5922), .Y(n2066));
   INVX1 U2240 ( .A(n5921), .Y(puf_3_wire_3));
   INVX1 U2241 ( .A(n5920), .Y(n2068));
   INVX1 U2242 ( .A(n5952), .Y(n2069));
   INVX1 U2243 ( .A(n5951), .Y(n2070));
   INVX1 U2244 ( .A(n5950), .Y(n2071));
   BUFX2 U2245 ( .A(k_data[23]), .Y(n2072));
   INVX1 U2246 ( .A(n5967), .Y(n2073));
   INVX1 U2247 ( .A(n5966), .Y(n2074));
   AND2X2 U2248 ( .A(n5968),  .B(n5969), .Y(n5967));
   INVX1 U2249 ( .A(n5978), .Y(n2075));
   INVX1 U2250 ( .A(n5977), .Y(n2076));
   INVX1 U2251 ( .A(n5976), .Y(n2077));
   INVX1 U2252 ( .A(n5995), .Y(n2078));
   INVX1 U2253 ( .A(n5994), .Y(n2079));
   INVX1 U2254 ( .A(n6017), .Y(n2080));
   INVX1 U2255 ( .A(n6016), .Y(n2081));
   INVX1 U2256 ( .A(n6015), .Y(n2082));
   INVX1 U2257 ( .A(n6042), .Y(n2083));
   INVX1 U2258 ( .A(n6041), .Y(n2084));
   INVX1 U2259 ( .A(n6040), .Y(n2085));
   BUFX2 U2260 ( .A(k_data[15]), .Y(n2086));
   INVX1 U2261 ( .A(n6063), .Y(n2087));
   INVX1 U2262 ( .A(n6062), .Y(n2088));
   INVX1 U2263 ( .A(n6077), .Y(n2089));
   INVX1 U2264 ( .A(n6076), .Y(n2090));
   INVX1 U2265 ( .A(n6075), .Y(n2091));
   AND2X2 U2266 ( .A(n6078),  .B(n6079), .Y(n6077));
   INVX1 U2267 ( .A(n6104), .Y(n2092));
   INVX1 U2268 ( .A(n6103), .Y(n2093));
   INVX1 U2269 ( .A(n6102), .Y(n2094));
   AND2X2 U2270 ( .A(n6105),  .B(n6106), .Y(n6104));
   INVX1 U2271 ( .A(n4655), .Y(n2095));
   INVX1 U2272 ( .A(n4654), .Y(n2096));
   OR2X2 U2273 ( .A(n4656),  .B(n4657), .Y(n4655));
   AND2X1 U2274 ( .A(n5805),  .B(n4705), .Y(n5846));
   INVX1 U2275 ( .A(n5846), .Y(n2097));
   AND2X1 U2276 ( .A(n5788),  .B(t_ctr_reg[5]), .Y(n6109));
   INVX1 U2277 ( .A(n6109), .Y(n2098));
   INVX1 U2278 ( .A(n6083), .Y(n2099));
   INVX1 U2279 ( .A(n6082), .Y(n2100));
   INVX1 U2280 ( .A(n5781), .Y(n2101));
   AND2X1 U2281 ( .A(n5859),  .B(n5917), .Y(n5781));
   BUFX2 U2282 ( .A(n4699), .Y(n2102));
   AND2X1 U2283 ( .A(n6001),  .B(n4711), .Y(n5886));
   INVX1 U2284 ( .A(n5886), .Y(n2103));
   AND2X1 U2285 ( .A(n6061),  .B(n6001), .Y(n5883));
   INVX1 U2286 ( .A(n5883), .Y(n2104));
   AND2X1 U2287 ( .A(n6001),  .B(n6000), .Y(n6068));
   INVX1 U2288 ( .A(n6068), .Y(n2105));
   AND2X1 U2289 ( .A(n6021),  .B(n4711), .Y(n5904));
   INVX1 U2290 ( .A(n5904), .Y(n2106));
   AND2X1 U2291 ( .A(n5885),  .B(n4711), .Y(n6038));
   INVX1 U2292 ( .A(n6038), .Y(n2107));
   INVX1 U2293 ( .A(n5926), .Y(n2108));
   AND2X1 U2294 ( .A(n2782),  .B(n2116), .Y(n5926));
   AND2X1 U2295 ( .A(n5807),  .B(n5789), .Y(n5779));
   INVX1 U2296 ( .A(n5779), .Y(n2109));
   AND2X1 U2297 ( .A(n2889),  .B(n2655), .Y(n5755));
   INVX1 U2298 ( .A(n5755), .Y(n2110));
   AND2X1 U2299 ( .A(n5860),  .B(n5763), .Y(n5838));
   INVX1 U2300 ( .A(n5838), .Y(n2111));
   AND2X1 U2301 ( .A(n5814),  .B(n5763), .Y(n5778));
   INVX1 U2302 ( .A(n5778), .Y(n2112));
   AND2X1 U2303 ( .A(n5998),  .B(n4711), .Y(n5914));
   INVX1 U2304 ( .A(n5914), .Y(n2113));
   INVX1 U2305 ( .A(n5769), .Y(n2114));
   AND2X1 U2306 ( .A(n5925),  .B(n4711), .Y(n5769));
   INVX1 U2307 ( .A(n5889), .Y(n2115));
   AND2X1 U2308 ( .A(n6109),  .B(n4705), .Y(n5889));
   AND2X1 U2309 ( .A(n5998),  .B(n4705), .Y(n5925));
   INVX1 U2310 ( .A(n5925), .Y(n2116));
   INVX1 U2311 ( .A(n4170), .Y(n2117));
   INVX1 U2312 ( .A(n4154), .Y(n2118));
   INVX1 U2313 ( .A(n2118), .Y(n2119));
   INVX1 U2314 ( .A(n4152), .Y(n2120));
   INVX1 U2315 ( .A(n2120), .Y(n2121));
   INVX1 U2316 ( .A(n4159), .Y(n2122));
   INVX1 U2317 ( .A(n2122), .Y(n2123));
   INVX1 U2318 ( .A(n4153), .Y(n2124));
   INVX1 U2319 ( .A(n2124), .Y(n2125));
   AND2X2 U2320 ( .A(n3041),  .B(n5676), .Y(n4718));
   INVX2 U2321 ( .A(n3088), .Y(puf_4_wire_3));
   INVX1 U2322 ( .A(n3116), .Y(n2127));
   AND2X1 U2323 ( .A(N686),  .B(n3087), .Y(n4925));
   INVX1 U2324 ( .A(n4925), .Y(n2128));
   AND2X1 U2325 ( .A(N698),  .B(n3087), .Y(n4949));
   INVX1 U2326 ( .A(n4949), .Y(n2129));
   AND2X1 U2327 ( .A(N715),  .B(n3086), .Y(n5047));
   INVX1 U2328 ( .A(n5047), .Y(n2130));
   AND2X1 U2329 ( .A(N731),  .B(n3087), .Y(n5079));
   INVX1 U2330 ( .A(n5079), .Y(n2131));
   AND2X1 U2331 ( .A(N771),  .B(n3086), .Y(n5223));
   INVX1 U2332 ( .A(n5223), .Y(n2132));
   AND2X1 U2333 ( .A(N553),  .B(n3087), .Y(n5427));
   INVX1 U2334 ( .A(n5427), .Y(n2133));
   AND2X1 U2335 ( .A(N583),  .B(n3086), .Y(n5551));
   INVX1 U2336 ( .A(n5551), .Y(n2134));
   BUFX2 U2337 ( .A(n4014), .Y(n2135));
   BUFX2 U2338 ( .A(n3630), .Y(n2136));
   BUFX2 U2339 ( .A(n3246), .Y(n2137));
   AND2X1 U2340 ( .A(N688),  .B(n3087), .Y(n4929));
   INVX1 U2341 ( .A(n4929), .Y(n2138));
   AND2X1 U2342 ( .A(N699),  .B(n3087), .Y(n4951));
   INVX1 U2343 ( .A(n4951), .Y(n2139));
   AND2X1 U2344 ( .A(N716),  .B(n3086), .Y(n5049));
   INVX1 U2345 ( .A(n5049), .Y(n2140));
   AND2X1 U2346 ( .A(N732),  .B(n3087), .Y(n5081));
   INVX1 U2347 ( .A(n5081), .Y(n2141));
   AND2X1 U2348 ( .A(N772),  .B(n3087), .Y(n5225));
   INVX1 U2349 ( .A(n5225), .Y(n2142));
   AND2X1 U2350 ( .A(N554),  .B(n3085), .Y(n5429));
   INVX1 U2351 ( .A(n5429), .Y(n2143));
   AND2X1 U2352 ( .A(N585),  .B(n3085), .Y(n5555));
   INVX1 U2353 ( .A(n5555), .Y(n2144));
   BUFX2 U2354 ( .A(n3886), .Y(n2145));
   BUFX2 U2355 ( .A(n3694), .Y(n2146));
   BUFX2 U2356 ( .A(n3310), .Y(n2147));
   BUFX2 U2357 ( .A(n3628), .Y(n2148));
   BUFX2 U2358 ( .A(n3244), .Y(n2149));
   BUFX2 U2359 ( .A(n4010), .Y(n2150));
   AND2X1 U2360 ( .A(N693),  .B(n3085), .Y(n4939));
   INVX1 U2361 ( .A(n4939), .Y(n2151));
   AND2X1 U2362 ( .A(N703),  .B(n3086), .Y(n4959));
   INVX1 U2363 ( .A(n4959), .Y(n2152));
   AND2X1 U2364 ( .A(N718),  .B(n3086), .Y(n5053));
   INVX1 U2365 ( .A(n5053), .Y(n2153));
   AND2X1 U2366 ( .A(N733),  .B(n3087), .Y(n5083));
   INVX1 U2367 ( .A(n5083), .Y(n2154));
   AND2X1 U2368 ( .A(N775),  .B(n3085), .Y(n5295));
   INVX1 U2369 ( .A(n5295), .Y(n2155));
   AND2X1 U2370 ( .A(N557),  .B(n3086), .Y(n5435));
   INVX1 U2371 ( .A(n5435), .Y(n2156));
   AND2X1 U2372 ( .A(N586),  .B(n3085), .Y(n5557));
   INVX1 U2373 ( .A(n5557), .Y(n2157));
   BUFX2 U2374 ( .A(n3822), .Y(n2158));
   BUFX2 U2375 ( .A(n3566), .Y(n2159));
   BUFX2 U2376 ( .A(n3884), .Y(n2160));
   BUFX2 U2377 ( .A(n3372), .Y(n2161));
   BUFX2 U2378 ( .A(n4008), .Y(n2162));
   BUFX2 U2379 ( .A(n3624), .Y(n2163));
   BUFX2 U2380 ( .A(n3240), .Y(n2164));
   BUFX2 U2381 ( .A(n4070), .Y(n2165));
   BUFX2 U2382 ( .A(n3686), .Y(n2166));
   BUFX2 U2383 ( .A(n3302), .Y(n2167));
   BUFX2 U2384 ( .A(n4911), .Y(n2168));
   BUFX2 U2385 ( .A(n5481), .Y(n2169));
   BUFX2 U2386 ( .A(n5593), .Y(n2170));
   AND2X1 U2387 ( .A(N700),  .B(n3087), .Y(n4953));
   INVX1 U2388 ( .A(n4953), .Y(n2171));
   AND2X1 U2389 ( .A(N719),  .B(n3086), .Y(n5055));
   INVX1 U2390 ( .A(n5055), .Y(n2172));
   AND2X1 U2391 ( .A(N736),  .B(n3087), .Y(n5089));
   INVX1 U2392 ( .A(n5089), .Y(n2173));
   AND2X1 U2393 ( .A(N776),  .B(n3087), .Y(n5297));
   INVX1 U2394 ( .A(n5297), .Y(n2174));
   AND2X1 U2395 ( .A(N558),  .B(n3086), .Y(n5437));
   INVX1 U2396 ( .A(n5437), .Y(n2175));
   AND2X1 U2397 ( .A(N594),  .B(n3086), .Y(n5573));
   INVX1 U2398 ( .A(n5573), .Y(n2176));
   BUFX2 U2399 ( .A(n3758), .Y(n2177));
   BUFX2 U2400 ( .A(n3374), .Y(n2178));
   BUFX2 U2401 ( .A(n3182), .Y(n2179));
   BUFX2 U2402 ( .A(n3820), .Y(n2180));
   BUFX2 U2403 ( .A(n3564), .Y(n2181));
   BUFX2 U2404 ( .A(n3308), .Y(n2182));
   BUFX2 U2405 ( .A(n4006), .Y(n2183));
   BUFX2 U2406 ( .A(n3878), .Y(n2184));
   BUFX2 U2407 ( .A(n3622), .Y(n2185));
   BUFX2 U2408 ( .A(n3238), .Y(n2186));
   BUFX2 U2409 ( .A(n4068), .Y(n2187));
   BUFX2 U2410 ( .A(n3684), .Y(n2188));
   BUFX2 U2411 ( .A(n4913), .Y(n2189));
   BUFX2 U2412 ( .A(n4969), .Y(n2190));
   BUFX2 U2413 ( .A(n5563), .Y(n2191));
   BUFX2 U2414 ( .A(n5603), .Y(n2192));
   AND2X1 U2415 ( .A(N701),  .B(n3085), .Y(n4955));
   INVX1 U2416 ( .A(n4955), .Y(n2193));
   AND2X1 U2417 ( .A(N739),  .B(n3087), .Y(n5095));
   INVX1 U2418 ( .A(n5095), .Y(n2194));
   AND2X1 U2419 ( .A(N779),  .B(n3085), .Y(n5303));
   INVX1 U2420 ( .A(n5303), .Y(n2195));
   AND2X1 U2421 ( .A(N561),  .B(n3087), .Y(n5443));
   INVX1 U2422 ( .A(n5443), .Y(n2196));
   AND2X1 U2423 ( .A(N596),  .B(n3086), .Y(n5577));
   INVX1 U2424 ( .A(n5577), .Y(n2197));
   AND2X1 U2425 ( .A(N648),  .B(n3086), .Y(n4785));
   INVX1 U2426 ( .A(n4785), .Y(n2198));
   BUFX2 U2427 ( .A(n4142), .Y(n2199));
   BUFX2 U2428 ( .A(n3756), .Y(n2200));
   BUFX2 U2429 ( .A(n3500), .Y(n2201));
   BUFX2 U2430 ( .A(n3180), .Y(n2202));
   BUFX2 U2431 ( .A(n3562), .Y(n2203));
   BUFX2 U2432 ( .A(n3370), .Y(n2204));
   BUFX2 U2433 ( .A(n3816), .Y(n2205));
   BUFX2 U2434 ( .A(n4004), .Y(n2206));
   BUFX2 U2435 ( .A(n3876), .Y(n2207));
   BUFX2 U2436 ( .A(n3620), .Y(n2208));
   BUFX2 U2437 ( .A(n3236), .Y(n2209));
   BUFX2 U2438 ( .A(n4066), .Y(n2210));
   BUFX2 U2439 ( .A(n3682), .Y(n2211));
   BUFX2 U2440 ( .A(n3298), .Y(n2212));
   BUFX2 U2441 ( .A(n3854), .Y(n2213));
   BUFX2 U2442 ( .A(n3278), .Y(n2214));
   BUFX2 U2443 ( .A(n4933), .Y(n2215));
   BUFX2 U2444 ( .A(n5041), .Y(n2216));
   BUFX2 U2445 ( .A(n5425), .Y(n2217));
   BUFX2 U2446 ( .A(n5567), .Y(n2218));
   BUFX2 U2447 ( .A(n5597), .Y(n2219));
   BUFX2 U2448 ( .A(n5704), .Y(n2220));
   AND2X1 U2449 ( .A(N704),  .B(n3085), .Y(n4961));
   INVX1 U2450 ( .A(n4961), .Y(n2221));
   AND2X1 U2451 ( .A(N727),  .B(n3085), .Y(n5071));
   INVX1 U2452 ( .A(n5071), .Y(n2222));
   AND2X1 U2453 ( .A(N740),  .B(n3087), .Y(n5097));
   INVX1 U2454 ( .A(n5097), .Y(n2223));
   AND2X1 U2455 ( .A(N790),  .B(n3086), .Y(n5325));
   INVX1 U2456 ( .A(n5325), .Y(n2224));
   AND2X1 U2457 ( .A(N570),  .B(n3085), .Y(n5461));
   INVX1 U2458 ( .A(n5461), .Y(n2225));
   AND2X1 U2459 ( .A(N601),  .B(n3086), .Y(n5587));
   INVX1 U2460 ( .A(n5587), .Y(n2226));
   AND2X1 U2461 ( .A(N630),  .B(n3085), .Y(n5710));
   INVX1 U2462 ( .A(n5710), .Y(n2227));
   AND2X1 U2463 ( .A(N652),  .B(n3086), .Y(n4793));
   INVX1 U2464 ( .A(n4793), .Y(n2228));
   BUFX2 U2465 ( .A(n4078), .Y(n2229));
   BUFX2 U2466 ( .A(n3438), .Y(n2230));
   BUFX2 U2467 ( .A(n4140), .Y(n2231));
   BUFX2 U2468 ( .A(n3692), .Y(n2232));
   BUFX2 U2469 ( .A(n3754), .Y(n2233));
   BUFX2 U2470 ( .A(n3944), .Y(n2234));
   BUFX2 U2471 ( .A(n3496), .Y(n2235));
   BUFX2 U2472 ( .A(n3368), .Y(n2236));
   BUFX2 U2473 ( .A(n3814), .Y(n2237));
   BUFX2 U2474 ( .A(n3300), .Y(n2238));
   BUFX2 U2475 ( .A(n4002), .Y(n2239));
   BUFX2 U2476 ( .A(n3874), .Y(n2240));
   BUFX2 U2477 ( .A(n3618), .Y(n2241));
   BUFX2 U2478 ( .A(n3234), .Y(n2242));
   BUFX2 U2479 ( .A(n4062), .Y(n2243));
   BUFX2 U2480 ( .A(n3676), .Y(n2244));
   BUFX2 U2481 ( .A(n3548), .Y(n2245));
   BUFX2 U2482 ( .A(n3420), .Y(n2246));
   BUFX2 U2483 ( .A(n3162), .Y(n2247));
   BUFX2 U2484 ( .A(n4114), .Y(n2248));
   BUFX2 U2485 ( .A(n3984), .Y(n2249));
   BUFX2 U2486 ( .A(n3728), .Y(n2250));
   BUFX2 U2487 ( .A(n3600), .Y(n2251));
   BUFX2 U2488 ( .A(n3790), .Y(n2252));
   BUFX2 U2489 ( .A(n3470), .Y(n2253));
   BUFX2 U2490 ( .A(n3342), .Y(n2254));
   BUFX2 U2491 ( .A(n3214), .Y(n2255));
   BUFX2 U2492 ( .A(n3916), .Y(n2256));
   BUFX2 U2493 ( .A(n4937), .Y(n2257));
   BUFX2 U2494 ( .A(n5197), .Y(n2258));
   BUFX2 U2495 ( .A(n5315), .Y(n2259));
   BUFX2 U2496 ( .A(n5431), .Y(n2260));
   BUFX2 U2497 ( .A(n5569), .Y(n2261));
   BUFX2 U2498 ( .A(n5702), .Y(n2262));
   BUFX2 U2499 ( .A(n4805), .Y(n2263));
   AND2X1 U2500 ( .A(N646),  .B(n3086), .Y(n4715));
   INVX1 U2501 ( .A(n4715), .Y(n2264));
   AND2X1 U2502 ( .A(N714),  .B(n3085), .Y(n5045));
   INVX1 U2503 ( .A(n5045), .Y(n2265));
   AND2X1 U2504 ( .A(N744),  .B(n3087), .Y(n5169));
   INVX1 U2505 ( .A(n5169), .Y(n2266));
   AND2X1 U2506 ( .A(N791),  .B(n3085), .Y(n5327));
   INVX1 U2507 ( .A(n5327), .Y(n2267));
   AND2X1 U2508 ( .A(N562),  .B(n3087), .Y(n5445));
   INVX1 U2509 ( .A(n5445), .Y(n2268));
   AND2X1 U2510 ( .A(N587),  .B(n3087), .Y(n5559));
   INVX1 U2511 ( .A(n5559), .Y(n2269));
   AND2X1 U2512 ( .A(N634),  .B(n3087), .Y(n5718));
   INVX1 U2513 ( .A(n5718), .Y(n2270));
   BUFX2 U2514 ( .A(n3502), .Y(n2271));
   BUFX2 U2515 ( .A(n4076), .Y(n2272));
   BUFX2 U2516 ( .A(n3436), .Y(n2273));
   BUFX2 U2517 ( .A(n4138), .Y(n2274));
   BUFX2 U2518 ( .A(n3178), .Y(n2275));
   BUFX2 U2519 ( .A(n3752), .Y(n2276));
   BUFX2 U2520 ( .A(n3560), .Y(n2277));
   BUFX2 U2521 ( .A(n3942), .Y(n2278));
   BUFX2 U2522 ( .A(n3494), .Y(n2279));
   BUFX2 U2523 ( .A(n3366), .Y(n2280));
   BUFX2 U2524 ( .A(n3812), .Y(n2281));
   BUFX2 U2525 ( .A(n4000), .Y(n2282));
   BUFX2 U2526 ( .A(n3872), .Y(n2283));
   BUFX2 U2527 ( .A(n3616), .Y(n2284));
   BUFX2 U2528 ( .A(n3232), .Y(n2285));
   BUFX2 U2529 ( .A(n3678), .Y(n2286));
   BUFX2 U2530 ( .A(n3294), .Y(puf_5_wire_3));
   BUFX2 U2531 ( .A(n4060), .Y(n2288));
   BUFX2 U2532 ( .A(n3542), .Y(n2289));
   BUFX2 U2533 ( .A(n3158), .Y(n2290));
   BUFX2 U2534 ( .A(n4110), .Y(n2291));
   BUFX2 U2535 ( .A(n3918), .Y(n2292));
   BUFX2 U2536 ( .A(n3662), .Y(n2293));
   BUFX2 U2537 ( .A(n3852), .Y(n2294));
   BUFX2 U2538 ( .A(n3724), .Y(n2295));
   BUFX2 U2539 ( .A(n3468), .Y(n2296));
   BUFX2 U2540 ( .A(n3276), .Y(n2297));
   BUFX2 U2541 ( .A(n3338), .Y(n2298));
   BUFX2 U2542 ( .A(n3974), .Y(n2299));
   BUFX2 U2543 ( .A(n3782), .Y(n2300));
   BUFX2 U2544 ( .A(n3590), .Y(n2301));
   BUFX2 U2545 ( .A(n3398), .Y(n2302));
   BUFX2 U2546 ( .A(n3206), .Y(n2303));
   BUFX2 U2547 ( .A(n4036), .Y(n2304));
   BUFX2 U2548 ( .A(n4915), .Y(n2305));
   BUFX2 U2549 ( .A(n4957), .Y(n2306));
   BUFX2 U2550 ( .A(n5091), .Y(n2307));
   BUFX2 U2551 ( .A(n5199), .Y(n2308));
   BUFX2 U2552 ( .A(n5321), .Y(n2309));
   BUFX2 U2553 ( .A(n5471), .Y(n2310));
   BUFX2 U2554 ( .A(n5571), .Y(n2311));
   BUFX2 U2555 ( .A(n5599), .Y(n2312));
   BUFX2 U2556 ( .A(n5706), .Y(n2313));
   BUFX2 U2557 ( .A(n4807), .Y(n2314));
   AND2X1 U2558 ( .A(N722),  .B(n3085), .Y(n5061));
   INVX1 U2559 ( .A(n5061), .Y(n2315));
   AND2X1 U2560 ( .A(N751),  .B(n3087), .Y(n5183));
   INVX1 U2561 ( .A(n5183), .Y(n2316));
   AND2X1 U2562 ( .A(N792),  .B(n3087), .Y(n5329));
   INVX1 U2563 ( .A(n5329), .Y(n2317));
   AND2X1 U2564 ( .A(N567),  .B(n3086), .Y(n5455));
   INVX1 U2565 ( .A(n5455), .Y(n2318));
   AND2X1 U2566 ( .A(N588),  .B(n3086), .Y(n5561));
   INVX1 U2567 ( .A(n5561), .Y(n2319));
   AND2X1 U2568 ( .A(N621),  .B(n3086), .Y(n5692));
   INVX1 U2569 ( .A(n5692), .Y(n2320));
   AND2X1 U2570 ( .A(N667),  .B(n3087), .Y(n4823));
   INVX1 U2571 ( .A(n4823), .Y(n2321));
   BUFX2 U2572 ( .A(n4012), .Y(n2322));
   BUFX2 U2573 ( .A(n3882), .Y(n2323));
   BUFX2 U2574 ( .A(n3626), .Y(n2324));
   BUFX2 U2575 ( .A(n3498), .Y(n2325));
   BUFX2 U2576 ( .A(n3242), .Y(n2326));
   BUFX2 U2577 ( .A(n4136), .Y(n2327));
   BUFX2 U2578 ( .A(n3750), .Y(n2328));
   BUFX2 U2579 ( .A(n3558), .Y(n2329));
   BUFX2 U2580 ( .A(n3940), .Y(n2330));
   BUFX2 U2581 ( .A(n3492), .Y(n2331));
   BUFX2 U2582 ( .A(n3364), .Y(n2332));
   BUFX2 U2583 ( .A(n4064), .Y(n2333));
   BUFX2 U2584 ( .A(n3680), .Y(n2334));
   BUFX2 U2585 ( .A(n3296), .Y(n2335));
   BUFX2 U2586 ( .A(n3998), .Y(n2336));
   BUFX2 U2587 ( .A(n3806), .Y(n2337));
   BUFX2 U2588 ( .A(n3614), .Y(n2338));
   BUFX2 U2589 ( .A(n3422), .Y(n2339));
   BUFX2 U2590 ( .A(n3230), .Y(n2340));
   BUFX2 U2591 ( .A(n3866), .Y(n2341));
   BUFX2 U2592 ( .A(n3160), .Y(n2342));
   BUFX2 U2593 ( .A(n3540), .Y(n2343));
   BUFX2 U2594 ( .A(n4112), .Y(n2344));
   BUFX2 U2595 ( .A(n4046), .Y(n2345));
   BUFX2 U2596 ( .A(n3726), .Y(n2346));
   BUFX2 U2597 ( .A(n3660), .Y(n2347));
   BUFX2 U2598 ( .A(n3340), .Y(n2348));
   BUFX2 U2599 ( .A(n3914), .Y(n2349));
   BUFX2 U2600 ( .A(n3466), .Y(n2350));
   BUFX2 U2601 ( .A(n3274), .Y(n2351));
   BUFX2 U2602 ( .A(n3972), .Y(n2352));
   BUFX2 U2603 ( .A(n3780), .Y(n2353));
   BUFX2 U2604 ( .A(n3588), .Y(n2354));
   BUFX2 U2605 ( .A(n3396), .Y(n2355));
   BUFX2 U2606 ( .A(n3204), .Y(n2356));
   BUFX2 U2607 ( .A(n3842), .Y(n2357));
   BUFX2 U2608 ( .A(n3136), .Y(n2358));
   BUFX2 U2609 ( .A(n4917), .Y(n2359));
   BUFX2 U2610 ( .A(n4965), .Y(n2360));
   BUFX2 U2611 ( .A(n5093), .Y(n2361));
   BUFX2 U2612 ( .A(n5211), .Y(n2362));
   BUFX2 U2613 ( .A(n5323), .Y(n2363));
   BUFX2 U2614 ( .A(n5475), .Y(n2364));
   BUFX2 U2615 ( .A(n5575), .Y(n2365));
   BUFX2 U2616 ( .A(n5605), .Y(n2366));
   BUFX2 U2617 ( .A(n5708), .Y(n2367));
   BUFX2 U2618 ( .A(n4809), .Y(n2368));
   AND2X1 U2619 ( .A(N720),  .B(n3086), .Y(n5057));
   INVX1 U2620 ( .A(n5057), .Y(n2369));
   AND2X1 U2621 ( .A(N752),  .B(n3087), .Y(n5185));
   INVX1 U2622 ( .A(n5185), .Y(n2370));
   AND2X1 U2623 ( .A(N780),  .B(n3086), .Y(n5305));
   INVX1 U2624 ( .A(n5305), .Y(n2371));
   AND2X1 U2625 ( .A(N568),  .B(n3087), .Y(n5457));
   INVX1 U2626 ( .A(n5457), .Y(n2372));
   AND2X1 U2627 ( .A(N590),  .B(n3087), .Y(n5565));
   INVX1 U2628 ( .A(n5565), .Y(n2373));
   AND2X1 U2629 ( .A(N624),  .B(n3085), .Y(n5698));
   INVX1 U2630 ( .A(n5698), .Y(n2374));
   AND2X1 U2631 ( .A(N653),  .B(n3086), .Y(n4795));
   INVX1 U2632 ( .A(n4795), .Y(n2375));
   AND2X1 U2633 ( .A(N669),  .B(n3085), .Y(n4827));
   INVX1 U2634 ( .A(n4827), .Y(n2376));
   BUFX2 U2635 ( .A(n4074), .Y(n2377));
   BUFX2 U2636 ( .A(n3818), .Y(n2378));
   BUFX2 U2637 ( .A(n3690), .Y(n2379));
   BUFX2 U2638 ( .A(n3434), .Y(n2380));
   BUFX2 U2639 ( .A(n3306), .Y(n2381));
   BUFX2 U2640 ( .A(n3176), .Y(n2382));
   BUFX2 U2641 ( .A(n4134), .Y(n2383));
   BUFX2 U2642 ( .A(n3748), .Y(n2384));
   BUFX2 U2643 ( .A(n3938), .Y(n2385));
   BUFX2 U2644 ( .A(n3490), .Y(n2386));
   BUFX2 U2645 ( .A(n3362), .Y(n2387));
   BUFX2 U2646 ( .A(n3870), .Y(n2388));
   BUFX2 U2647 ( .A(n3996), .Y(n2389));
   BUFX2 U2648 ( .A(n3804), .Y(n2390));
   BUFX2 U2649 ( .A(n3612), .Y(n2391));
   BUFX2 U2650 ( .A(n3228), .Y(n2392));
   BUFX2 U2651 ( .A(n4058), .Y(n2393));
   BUFX2 U2652 ( .A(n3674), .Y(n2394));
   BUFX2 U2653 ( .A(n3546), .Y(n2395));
   BUFX2 U2654 ( .A(n3418), .Y(n2396));
   BUFX2 U2655 ( .A(n3290), .Y(n2397));
   BUFX2 U2656 ( .A(n3156), .Y(n2398));
   BUFX2 U2657 ( .A(n4108), .Y(n2399));
   BUFX2 U2658 ( .A(n3850), .Y(n2400));
   BUFX2 U2659 ( .A(n3722), .Y(n2401));
   BUFX2 U2660 ( .A(n3912), .Y(n2402));
   BUFX2 U2661 ( .A(n3464), .Y(n2403));
   BUFX2 U2662 ( .A(n3336), .Y(n2404));
   BUFX2 U2663 ( .A(n3970), .Y(n2405));
   BUFX2 U2664 ( .A(n3778), .Y(n2406));
   BUFX2 U2665 ( .A(n3650), .Y(n2407));
   BUFX2 U2666 ( .A(n3522), .Y(n2408));
   BUFX2 U2667 ( .A(n3394), .Y(n2409));
   BUFX2 U2668 ( .A(n3202), .Y(n2410));
   BUFX2 U2669 ( .A(n4032), .Y(n2411));
   BUFX2 U2670 ( .A(n3584), .Y(n2412));
   BUFX2 U2671 ( .A(n3264), .Y(n2413));
   BUFX2 U2672 ( .A(n3134), .Y(n2414));
   BUFX2 U2673 ( .A(n4919), .Y(n2415));
   BUFX2 U2674 ( .A(n5043), .Y(n2416));
   BUFX2 U2675 ( .A(n5167), .Y(n2417));
   BUFX2 U2676 ( .A(n5213), .Y(n2418));
   BUFX2 U2677 ( .A(n5335), .Y(n2419));
   BUFX2 U2678 ( .A(n5479), .Y(n2420));
   BUFX2 U2679 ( .A(n5581), .Y(n2421));
   BUFX2 U2680 ( .A(n5712), .Y(n2422));
   BUFX2 U2681 ( .A(n4811), .Y(n2423));
   BUFX2 U2682 ( .A(n5827), .Y(n2424));
   AND2X1 U2683 ( .A(N705),  .B(n3086), .Y(n4963));
   INVX1 U2684 ( .A(n4963), .Y(n2425));
   AND2X1 U2685 ( .A(N725),  .B(n3086), .Y(n5067));
   INVX1 U2686 ( .A(n5067), .Y(n2426));
   AND2X1 U2687 ( .A(N755),  .B(n3087), .Y(n5191));
   INVX1 U2688 ( .A(n5191), .Y(n2427));
   AND2X1 U2689 ( .A(N781),  .B(n3085), .Y(n5307));
   INVX1 U2690 ( .A(n5307), .Y(n2428));
   AND2X1 U2691 ( .A(N571),  .B(n3085), .Y(n5463));
   INVX1 U2692 ( .A(n5463), .Y(n2429));
   AND2X1 U2693 ( .A(N602),  .B(n3085), .Y(n5589));
   INVX1 U2694 ( .A(n5589), .Y(n2430));
   AND2X1 U2695 ( .A(N637),  .B(n3086), .Y(n5724));
   INVX1 U2696 ( .A(n5724), .Y(n2431));
   AND2X1 U2697 ( .A(N671),  .B(n3086), .Y(n4831));
   INVX1 U2698 ( .A(n4831), .Y(n2432));
   BUFX2 U2699 ( .A(n4072), .Y(n2433));
   BUFX2 U2700 ( .A(n3880), .Y(n2434));
   BUFX2 U2701 ( .A(n3688), .Y(n2435));
   BUFX2 U2702 ( .A(n3432), .Y(n2436));
   BUFX2 U2703 ( .A(n3304), .Y(n2437));
   BUFX2 U2704 ( .A(n3174), .Y(n2438));
   BUFX2 U2705 ( .A(n4132), .Y(n2439));
   BUFX2 U2706 ( .A(n3746), .Y(n2440));
   BUFX2 U2707 ( .A(n3936), .Y(n2441));
   BUFX2 U2708 ( .A(n3488), .Y(n2442));
   BUFX2 U2709 ( .A(n3360), .Y(n2443));
   BUFX2 U2710 ( .A(n3994), .Y(n2444));
   BUFX2 U2711 ( .A(n3802), .Y(n2445));
   BUFX2 U2712 ( .A(n3610), .Y(n2446));
   BUFX2 U2713 ( .A(n3226), .Y(n2447));
   BUFX2 U2714 ( .A(n3864), .Y(n2448));
   BUFX2 U2715 ( .A(n3672), .Y(n2449));
   BUFX2 U2716 ( .A(n3544), .Y(n2450));
   BUFX2 U2717 ( .A(n3416), .Y(n2451));
   BUFX2 U2718 ( .A(n3288), .Y(n2452));
   BUFX2 U2719 ( .A(n4054), .Y(n2453));
   BUFX2 U2720 ( .A(n3154), .Y(n2454));
   BUFX2 U2721 ( .A(n4106), .Y(n2455));
   BUFX2 U2722 ( .A(n3720), .Y(n2456));
   BUFX2 U2723 ( .A(n3910), .Y(n2457));
   BUFX2 U2724 ( .A(n3462), .Y(n2458));
   BUFX2 U2725 ( .A(n3334), .Y(n2459));
   BUFX2 U2726 ( .A(n4034), .Y(n2460));
   BUFX2 U2727 ( .A(n3586), .Y(n2461));
   BUFX2 U2728 ( .A(n3266), .Y(n2462));
   BUFX2 U2729 ( .A(n3968), .Y(n2463));
   BUFX2 U2730 ( .A(n3776), .Y(n2464));
   BUFX2 U2731 ( .A(n3648), .Y(n2465));
   BUFX2 U2732 ( .A(n3520), .Y(n2466));
   BUFX2 U2733 ( .A(n3392), .Y(n2467));
   BUFX2 U2734 ( .A(n3200), .Y(n2468));
   BUFX2 U2735 ( .A(n3838), .Y(n2469));
   BUFX2 U2736 ( .A(n3132), .Y(n2470));
   BUFX2 U2737 ( .A(n5069), .Y(n2471));
   BUFX2 U2738 ( .A(n5171), .Y(n2472));
   BUFX2 U2739 ( .A(n5215), .Y(n2473));
   BUFX2 U2740 ( .A(n5337), .Y(n2474));
   BUFX2 U2741 ( .A(n5433), .Y(n2475));
   BUFX2 U2742 ( .A(n5680), .Y(n2476));
   BUFX2 U2743 ( .A(n5732), .Y(n2477));
   BUFX2 U2744 ( .A(n4813), .Y(n2478));
   BUFX2 U2745 ( .A(n5963), .Y(n2479));
   BUFX2 U2746 ( .A(k_data[26]), .Y(n2480));
   BUFX2 U2747 ( .A(n5928), .Y(n2481));
   AND2X2 U2748 ( .A(n5931),  .B(n5932), .Y(n5930));
   AND2X1 U2749 ( .A(N707),  .B(n3086), .Y(n4967));
   INVX1 U2750 ( .A(n4967), .Y(n2482));
   AND2X1 U2751 ( .A(N760),  .B(n3087), .Y(n5201));
   INVX1 U2752 ( .A(n5201), .Y(n2483));
   AND2X1 U2753 ( .A(N783),  .B(n3087), .Y(n5311));
   INVX1 U2754 ( .A(n5311), .Y(n2484));
   AND2X1 U2755 ( .A(N572),  .B(n3085), .Y(n5465));
   INVX1 U2756 ( .A(n5465), .Y(n2485));
   AND2X1 U2757 ( .A(N605),  .B(n3087), .Y(n5595));
   INVX1 U2758 ( .A(n5595), .Y(n2486));
   AND2X1 U2759 ( .A(N625),  .B(n3085), .Y(n5700));
   INVX1 U2760 ( .A(n5700), .Y(n2487));
   AND2X1 U2761 ( .A(N673),  .B(n3085), .Y(n4835));
   INVX1 U2762 ( .A(n4835), .Y(n2488));
   BUFX2 U2763 ( .A(n3430), .Y(n2489));
   BUFX2 U2764 ( .A(n3556), .Y(n2490));
   BUFX2 U2765 ( .A(n3172), .Y(n2491));
   BUFX2 U2766 ( .A(n4130), .Y(n2492));
   BUFX2 U2767 ( .A(n3744), .Y(n2493));
   BUFX2 U2768 ( .A(n3934), .Y(n2494));
   BUFX2 U2769 ( .A(n3486), .Y(n2495));
   BUFX2 U2770 ( .A(n3358), .Y(n2496));
   BUFX2 U2771 ( .A(n4056), .Y(n2497));
   BUFX2 U2772 ( .A(n3800), .Y(n2498));
   BUFX2 U2773 ( .A(n3608), .Y(n2499));
   BUFX2 U2774 ( .A(n3224), .Y(n2500));
   BUFX2 U2775 ( .A(n3990), .Y(n2501));
   BUFX2 U2776 ( .A(n3862), .Y(n2502));
   BUFX2 U2777 ( .A(n3670), .Y(n2503));
   BUFX2 U2778 ( .A(n3414), .Y(n2504));
   BUFX2 U2779 ( .A(n3286), .Y(n2505));
   BUFX2 U2780 ( .A(n3538), .Y(n2506));
   BUFX2 U2781 ( .A(n3152), .Y(n2507));
   BUFX2 U2782 ( .A(n3460), .Y(n2508));
   BUFX2 U2783 ( .A(n3840), .Y(n2509));
   BUFX2 U2784 ( .A(n4094), .Y(n2510));
   BUFX2 U2785 ( .A(n3966), .Y(n2511));
   BUFX2 U2786 ( .A(n3774), .Y(n2512));
   BUFX2 U2787 ( .A(n3646), .Y(n2513));
   BUFX2 U2788 ( .A(n3518), .Y(n2514));
   BUFX2 U2789 ( .A(n3326), .Y(n2515));
   BUFX2 U2790 ( .A(n3198), .Y(n2516));
   BUFX2 U2791 ( .A(n4028), .Y(n2517));
   BUFX2 U2792 ( .A(n3900), .Y(n2518));
   BUFX2 U2793 ( .A(n3708), .Y(n2519));
   BUFX2 U2794 ( .A(n3580), .Y(n2520));
   BUFX2 U2795 ( .A(n3388), .Y(n2521));
   BUFX2 U2796 ( .A(n3260), .Y(n2522));
   BUFX2 U2797 ( .A(n3130), .Y(n2523));
   BUFX2 U2798 ( .A(n4921), .Y(n2524));
   BUFX2 U2799 ( .A(n5051), .Y(n2525));
   BUFX2 U2800 ( .A(n5175), .Y(n2526));
   BUFX2 U2801 ( .A(n5217), .Y(n2527));
   BUFX2 U2802 ( .A(n5339), .Y(n2528));
   BUFX2 U2803 ( .A(n5447), .Y(n2529));
   BUFX2 U2804 ( .A(n5553), .Y(n2530));
   BUFX2 U2805 ( .A(n5714), .Y(n2531));
   BUFX2 U2806 ( .A(n4787), .Y(n2532));
   BUFX2 U2807 ( .A(n4815), .Y(n2533));
   BUFX2 U2808 ( .A(n5990), .Y(n2534));
   AND2X1 U2809 ( .A(n5855),  .B(n5856), .Y(n5852));
   INVX1 U2810 ( .A(n5852), .Y(n2535));
   AND2X1 U2811 ( .A(n5859),  .B(n4705), .Y(n6061));
   INVX1 U2812 ( .A(n6061), .Y(n2536));
   BUFX2 U2813 ( .A(k_data[25]), .Y(n2537));
   BUFX2 U2814 ( .A(n5940), .Y(n2538));
   AND2X2 U2815 ( .A(n5943),  .B(n5944), .Y(n5942));
   AND2X1 U2816 ( .A(N710),  .B(n3087), .Y(n5037));
   INVX1 U2817 ( .A(n5037), .Y(n2539));
   AND2X1 U2818 ( .A(N729),  .B(n3086), .Y(n5075));
   INVX1 U2819 ( .A(n5075), .Y(n2540));
   AND2X1 U2820 ( .A(N761),  .B(n3087), .Y(n5203));
   INVX1 U2821 ( .A(n5203), .Y(n2541));
   AND2X1 U2822 ( .A(N786),  .B(n3087), .Y(n5317));
   INVX1 U2823 ( .A(n5317), .Y(n2542));
   AND2X1 U2824 ( .A(N573),  .B(n3086), .Y(n5467));
   INVX1 U2825 ( .A(n5467), .Y(n2543));
   AND2X1 U2826 ( .A(N617),  .B(n3085), .Y(n5684));
   INVX1 U2827 ( .A(n5684), .Y(n2544));
   AND2X1 U2828 ( .A(N638),  .B(n3087), .Y(n5726));
   INVX1 U2829 ( .A(n5726), .Y(n2545));
   AND2X1 U2830 ( .A(N676),  .B(n3086), .Y(n4841));
   INVX1 U2831 ( .A(n4841), .Y(n2546));
   BUFX2 U2832 ( .A(n3428), .Y(n2547));
   BUFX2 U2833 ( .A(n3810), .Y(n2548));
   BUFX2 U2834 ( .A(n3554), .Y(n2549));
   BUFX2 U2835 ( .A(n3170), .Y(n2550));
   BUFX2 U2836 ( .A(n3484), .Y(n2551));
   BUFX2 U2837 ( .A(n3992), .Y(n2552));
   BUFX2 U2838 ( .A(n3926), .Y(n2553));
   BUFX2 U2839 ( .A(n3734), .Y(n2554));
   BUFX2 U2840 ( .A(n3606), .Y(n2555));
   BUFX2 U2841 ( .A(n3350), .Y(n2556));
   BUFX2 U2842 ( .A(n3222), .Y(n2557));
   BUFX2 U2843 ( .A(n4116), .Y(n2558));
   BUFX2 U2844 ( .A(n3860), .Y(n2559));
   BUFX2 U2845 ( .A(n3668), .Y(n2560));
   BUFX2 U2846 ( .A(n3412), .Y(n2561));
   BUFX2 U2847 ( .A(n3284), .Y(n2562));
   BUFX2 U2848 ( .A(n4050), .Y(n2563));
   BUFX2 U2849 ( .A(n3536), .Y(n2564));
   BUFX2 U2850 ( .A(n3150), .Y(n2565));
   BUFX2 U2851 ( .A(n3788), .Y(n2566));
   BUFX2 U2852 ( .A(n3458), .Y(n2567));
   BUFX2 U2853 ( .A(n4030), .Y(n2568));
   BUFX2 U2854 ( .A(n3902), .Y(n2569));
   BUFX2 U2855 ( .A(n3710), .Y(n2570));
   BUFX2 U2856 ( .A(n3582), .Y(n2571));
   BUFX2 U2857 ( .A(n3390), .Y(n2572));
   BUFX2 U2858 ( .A(n3262), .Y(n2573));
   BUFX2 U2859 ( .A(n4092), .Y(n2574));
   BUFX2 U2860 ( .A(n3964), .Y(n2575));
   BUFX2 U2861 ( .A(n3836), .Y(n2576));
   BUFX2 U2862 ( .A(n3644), .Y(n2577));
   BUFX2 U2863 ( .A(n3516), .Y(n2578));
   BUFX2 U2864 ( .A(n3324), .Y(n2579));
   BUFX2 U2865 ( .A(n3196), .Y(n2580));
   BUFX2 U2866 ( .A(n3768), .Y(n2581));
   BUFX2 U2867 ( .A(n4927), .Y(n2582));
   BUFX2 U2868 ( .A(n5059), .Y(n2583));
   BUFX2 U2869 ( .A(n5179), .Y(n2584));
   BUFX2 U2870 ( .A(n5219), .Y(n2585));
   BUFX2 U2871 ( .A(n5341), .Y(n2586));
   BUFX2 U2872 ( .A(n5449), .Y(n2587));
   BUFX2 U2873 ( .A(n5607), .Y(n2588));
   BUFX2 U2874 ( .A(n5734), .Y(n2589));
   BUFX2 U2875 ( .A(n4817), .Y(n2590));
   AND2X1 U2876 ( .A(t_ctr_reg[4]),  .B(n2715), .Y(n6074));
   INVX1 U2877 ( .A(n6074), .Y(n2591));
   AND2X1 U2878 ( .A(n5861),  .B(n2657), .Y(n5899));
   INVX1 U2879 ( .A(n5899), .Y(n2592));
   AND2X1 U2880 ( .A(n6021),  .B(t_ctr_reg[5]), .Y(n5807));
   INVX1 U2881 ( .A(n5807), .Y(n2593));
   AND2X1 U2882 ( .A(n4707),  .B(n4711), .Y(n5859));
   INVX1 U2883 ( .A(n5859), .Y(n2594));
   AND2X1 U2884 ( .A(n5885),  .B(t_ctr_reg[2]), .Y(n5936));
   INVX1 U2885 ( .A(n5936), .Y(n2595));
   AND2X1 U2886 ( .A(N711),  .B(n3086), .Y(n5039));
   INVX1 U2887 ( .A(n5039), .Y(n2596));
   AND2X1 U2888 ( .A(N746),  .B(n3087), .Y(n5173));
   INVX1 U2889 ( .A(n5173), .Y(n2597));
   AND2X1 U2890 ( .A(N793),  .B(n3085), .Y(n5331));
   INVX1 U2891 ( .A(n5331), .Y(n2598));
   AND2X1 U2892 ( .A(N574),  .B(n3087), .Y(n5469));
   INVX1 U2893 ( .A(n5469), .Y(n2599));
   AND2X1 U2894 ( .A(N608),  .B(n3086), .Y(n5601));
   INVX1 U2895 ( .A(n5601), .Y(n2600));
   AND2X1 U2896 ( .A(N674),  .B(n3085), .Y(n4837));
   INVX1 U2897 ( .A(n4837), .Y(n2601));
   BUFX2 U2898 ( .A(n3950), .Y(n2602));
   BUFX2 U2899 ( .A(n3426), .Y(n2603));
   BUFX2 U2900 ( .A(n3552), .Y(n2604));
   BUFX2 U2901 ( .A(n3168), .Y(n2605));
   BUFX2 U2902 ( .A(n3482), .Y(n2606));
   BUFX2 U2903 ( .A(n4118), .Y(n2607));
   BUFX2 U2904 ( .A(n3798), .Y(n2608));
   BUFX2 U2905 ( .A(n4052), .Y(n2609));
   BUFX2 U2906 ( .A(n3924), .Y(n2610));
   BUFX2 U2907 ( .A(n3732), .Y(n2611));
   BUFX2 U2908 ( .A(n3604), .Y(n2612));
   BUFX2 U2909 ( .A(n3348), .Y(n2613));
   BUFX2 U2910 ( .A(n3220), .Y(n2614));
   BUFX2 U2911 ( .A(n3986), .Y(n2615));
   BUFX2 U2912 ( .A(n3858), .Y(n2616));
   BUFX2 U2913 ( .A(n3666), .Y(n2617));
   BUFX2 U2914 ( .A(n3410), .Y(n2618));
   BUFX2 U2915 ( .A(n3282), .Y(n2619));
   BUFX2 U2916 ( .A(n3534), .Y(n2620));
   BUFX2 U2917 ( .A(n3148), .Y(n2621));
   BUFX2 U2918 ( .A(n3456), .Y(n2622));
   BUFX2 U2919 ( .A(n3772), .Y(n2623));
   BUFX2 U2920 ( .A(n4090), .Y(n2624));
   BUFX2 U2921 ( .A(n3962), .Y(n2625));
   BUFX2 U2922 ( .A(n3834), .Y(n2626));
   BUFX2 U2923 ( .A(n3642), .Y(n2627));
   BUFX2 U2924 ( .A(n3514), .Y(n2628));
   BUFX2 U2925 ( .A(n3322), .Y(n2629));
   BUFX2 U2926 ( .A(n3194), .Y(n2630));
   BUFX2 U2927 ( .A(n4024), .Y(n2631));
   BUFX2 U2928 ( .A(n3896), .Y(n2632));
   BUFX2 U2929 ( .A(n3704), .Y(n2633));
   BUFX2 U2930 ( .A(n3576), .Y(n2634));
   BUFX2 U2931 ( .A(n3384), .Y(n2635));
   BUFX2 U2932 ( .A(n3256), .Y(n2636));
   BUFX2 U2933 ( .A(n3128), .Y(n2637));
   AND2X1 U2934 ( .A(w_mem_inst_N713),  .B(n3094), .Y(n3112));
   INVX1 U2935 ( .A(n3112), .Y(n2638));
   BUFX2 U2936 ( .A(n4943), .Y(n2639));
   BUFX2 U2937 ( .A(n5063), .Y(n2640));
   BUFX2 U2938 ( .A(n5181), .Y(n2641));
   BUFX2 U2939 ( .A(n5221), .Y(n2642));
   BUFX2 U2940 ( .A(n5349), .Y(n2643));
   BUFX2 U2941 ( .A(n5451), .Y(n2644));
   BUFX2 U2942 ( .A(n5686), .Y(n2645));
   BUFX2 U2943 ( .A(n5716), .Y(n2646));
   BUFX2 U2944 ( .A(n4782), .Y(n2647));
   BUFX2 U2945 ( .A(n4819), .Y(n2648));
   BUFX2 U2946 ( .A(k_data[20]), .Y(n2649));
   BUFX2 U2947 ( .A(n5985), .Y(n2650));
   AND2X2 U2948 ( .A(n5988),  .B(n5989), .Y(n5987));
   AND2X1 U2949 ( .A(n6109),  .B(t_ctr_reg[3]), .Y(n5822));
   INVX1 U2950 ( .A(n5822), .Y(n2651));
   AND2X1 U2951 ( .A(n2954),  .B(n2781), .Y(n5792));
   INVX1 U2952 ( .A(n5792), .Y(n2652));
   AND2X1 U2953 ( .A(n5771),  .B(n2784), .Y(n5819));
   INVX1 U2954 ( .A(n5819), .Y(n2653));
   AND2X1 U2955 ( .A(n6021),  .B(t_ctr_reg[4]), .Y(n5860));
   INVX1 U2956 ( .A(n5860), .Y(n2654));
   AND2X1 U2957 ( .A(n5859),  .B(n4703), .Y(n5875));
   INVX1 U2958 ( .A(n5875), .Y(n2655));
   AND2X1 U2959 ( .A(n5786),  .B(n2849), .Y(n5754));
   INVX1 U2960 ( .A(n5754), .Y(n2656));
   AND2X1 U2961 ( .A(t_ctr_reg[1]),  .B(t_ctr_reg[0]), .Y(n6001));
   INVX1 U2962 ( .A(n6001), .Y(n2657));
   AND2X1 U2963 ( .A(N730),  .B(n3087), .Y(n5077));
   INVX1 U2964 ( .A(n5077), .Y(n2658));
   AND2X1 U2965 ( .A(N762),  .B(n3087), .Y(n5205));
   INVX1 U2966 ( .A(n5205), .Y(n2659));
   AND2X1 U2967 ( .A(N787),  .B(n3087), .Y(n5319));
   INVX1 U2968 ( .A(n5319), .Y(n2660));
   AND2X1 U2969 ( .A(N576),  .B(n3085), .Y(n5473));
   INVX1 U2970 ( .A(n5473), .Y(n2661));
   AND2X1 U2971 ( .A(N612),  .B(n3085), .Y(n5609));
   INVX1 U2972 ( .A(n5609), .Y(n2662));
   AND2X1 U2973 ( .A(N655),  .B(n3085), .Y(n4799));
   INVX1 U2974 ( .A(n4799), .Y(n2663));
   BUFX2 U2975 ( .A(n3948), .Y(n2664));
   BUFX2 U2976 ( .A(n4128), .Y(n2665));
   BUFX2 U2977 ( .A(n3808), .Y(n2666));
   BUFX2 U2978 ( .A(n3424), .Y(n2667));
   BUFX2 U2979 ( .A(n3550), .Y(n2668));
   BUFX2 U2980 ( .A(n3166), .Y(n2669));
   BUFX2 U2981 ( .A(n3480), .Y(n2670));
   BUFX2 U2982 ( .A(n3988), .Y(n2671));
   BUFX2 U2983 ( .A(n3922), .Y(n2672));
   BUFX2 U2984 ( .A(n3730), .Y(n2673));
   BUFX2 U2985 ( .A(n3602), .Y(n2674));
   BUFX2 U2986 ( .A(n3346), .Y(n2675));
   BUFX2 U2987 ( .A(n3218), .Y(n2676));
   BUFX2 U2988 ( .A(n4048), .Y(n2677));
   BUFX2 U2989 ( .A(n3856), .Y(n2678));
   BUFX2 U2990 ( .A(n3664), .Y(n2679));
   BUFX2 U2991 ( .A(n3408), .Y(n2680));
   BUFX2 U2992 ( .A(n3280), .Y(n2681));
   BUFX2 U2993 ( .A(n3532), .Y(n2682));
   BUFX2 U2994 ( .A(n3786), .Y(n2683));
   BUFX2 U2995 ( .A(n3146), .Y(n2684));
   BUFX2 U2996 ( .A(n4104), .Y(n2685));
   BUFX2 U2997 ( .A(n3454), .Y(n2686));
   BUFX2 U2998 ( .A(n4026), .Y(n2687));
   BUFX2 U2999 ( .A(n3898), .Y(puf_6_wire_3));
   BUFX2 U3000 ( .A(n3706), .Y(n2689));
   BUFX2 U3001 ( .A(n3578), .Y(n2690));
   BUFX2 U3002 ( .A(n3386), .Y(n2691));
   BUFX2 U3003 ( .A(n3258), .Y(n2692));
   BUFX2 U3004 ( .A(n4088), .Y(n2693));
   BUFX2 U3005 ( .A(n3960), .Y(n2694));
   BUFX2 U3006 ( .A(n3832), .Y(n2695));
   BUFX2 U3007 ( .A(n3640), .Y(n2696));
   BUFX2 U3008 ( .A(n3512), .Y(n2697));
   BUFX2 U3009 ( .A(n3320), .Y(n2698));
   BUFX2 U3010 ( .A(n3192), .Y(n2699));
   BUFX2 U3011 ( .A(n3766), .Y(n2700));
   AND2X1 U3012 ( .A(w_mem_inst_N712),  .B(n3094), .Y(n3110));
   INVX1 U3013 ( .A(n3110), .Y(n2701));
   BUFX2 U3014 ( .A(n5065), .Y(n2702));
   BUFX2 U3015 ( .A(n5187), .Y(n2703));
   BUFX2 U3016 ( .A(n5299), .Y(n2704));
   BUFX2 U3017 ( .A(n5343), .Y(n2705));
   BUFX2 U3018 ( .A(n5439), .Y(n2706));
   BUFX2 U3019 ( .A(n5579), .Y(n2707));
   BUFX2 U3020 ( .A(n5688), .Y(n2708));
   BUFX2 U3021 ( .A(n5722), .Y(n2709));
   BUFX2 U3022 ( .A(n4789), .Y(n2710));
   BUFX2 U3023 ( .A(n4825), .Y(n2711));
   AND2X1 U3024 ( .A(n6002),  .B(n4707), .Y(n5840));
   INVX1 U3025 ( .A(n5840), .Y(n2712));
   AND2X1 U3026 ( .A(n2889),  .B(n2781), .Y(n5903));
   INVX1 U3027 ( .A(n5903), .Y(n2713));
   AND2X1 U3028 ( .A(n5934),  .B(n4711), .Y(n5972));
   INVX1 U3029 ( .A(n5972), .Y(n2714));
   AND2X1 U3030 ( .A(t_ctr_reg[3]),  .B(n4703), .Y(n6021));
   INVX1 U3031 ( .A(n6021), .Y(n2715));
   INVX1 U3032 ( .A(n5849), .Y(n2716));
   AND2X1 U3033 ( .A(n2954),  .B(n2892), .Y(n5757));
   INVX1 U3034 ( .A(n5757), .Y(n2717));
   AND2X1 U3035 ( .A(n6117),  .B(t_ctr_reg[5]), .Y(n5821));
   INVX1 U3036 ( .A(n5821), .Y(n2718));
   AND2X1 U3037 ( .A(n2849),  .B(n2891), .Y(n5916));
   INVX1 U3038 ( .A(n5916), .Y(n2719));
   AND2X1 U3039 ( .A(t_ctr_reg[0]),  .B(n4701), .Y(n5763));
   INVX1 U3040 ( .A(n5763), .Y(n2720));
   AND2X1 U3041 ( .A(N689),  .B(n3087), .Y(n4931));
   INVX1 U3042 ( .A(n4931), .Y(n2721));
   AND2X1 U3043 ( .A(N763),  .B(n3087), .Y(n5207));
   INVX1 U3044 ( .A(n5207), .Y(n2722));
   AND2X1 U3045 ( .A(N794),  .B(n3087), .Y(n5333));
   INVX1 U3046 ( .A(n5333), .Y(n2723));
   AND2X1 U3047 ( .A(N578),  .B(n3086), .Y(n5477));
   INVX1 U3048 ( .A(n5477), .Y(n2724));
   AND2X1 U3049 ( .A(N614),  .B(n3086), .Y(n5678));
   INVX1 U3050 ( .A(n5678), .Y(n2725));
   AND2X1 U3051 ( .A(N657),  .B(n3087), .Y(n4803));
   INVX1 U3052 ( .A(n4803), .Y(n2726));
   BUFX2 U3053 ( .A(n3946), .Y(n2727));
   BUFX2 U3054 ( .A(n4126), .Y(n2728));
   BUFX2 U3055 ( .A(n3742), .Y(n2729));
   BUFX2 U3056 ( .A(n3868), .Y(n2730));
   BUFX2 U3057 ( .A(n3356), .Y(n2731));
   BUFX2 U3058 ( .A(n3478), .Y(n2732));
   BUFX2 U3059 ( .A(n3796), .Y(n2733));
   BUFX2 U3060 ( .A(n3920), .Y(n2734));
   BUFX2 U3061 ( .A(n3982), .Y(n2735));
   BUFX2 U3062 ( .A(n3598), .Y(n2736));
   BUFX2 U3063 ( .A(n3406), .Y(n2737));
   BUFX2 U3064 ( .A(n4044), .Y(n2738));
   BUFX2 U3065 ( .A(n3212), .Y(n2739));
   BUFX2 U3066 ( .A(n3658), .Y(n2740));
   BUFX2 U3067 ( .A(n3530), .Y(n2741));
   BUFX2 U3068 ( .A(n3272), .Y(n2742));
   BUFX2 U3069 ( .A(n3144), .Y(n2743));
   BUFX2 U3070 ( .A(n4102), .Y(n2744));
   BUFX2 U3071 ( .A(n3718), .Y(n2745));
   BUFX2 U3072 ( .A(n3332), .Y(n2746));
   BUFX2 U3073 ( .A(n3452), .Y(n2747));
   BUFX2 U3074 ( .A(n3770), .Y(n2748));
   BUFX2 U3075 ( .A(n4022), .Y(n2749));
   BUFX2 U3076 ( .A(n3894), .Y(n2750));
   BUFX2 U3077 ( .A(n3638), .Y(n2751));
   BUFX2 U3078 ( .A(n3510), .Y(n2752));
   BUFX2 U3079 ( .A(n3382), .Y(n2753));
   BUFX2 U3080 ( .A(n3254), .Y(n2754));
   BUFX2 U3081 ( .A(n3126), .Y(n2755));
   BUFX2 U3082 ( .A(n4084), .Y(n2756));
   BUFX2 U3083 ( .A(n3956), .Y(n2757));
   BUFX2 U3084 ( .A(n3828), .Y(n2758));
   BUFX2 U3085 ( .A(n3700), .Y(n2759));
   BUFX2 U3086 ( .A(n3572), .Y(n2760));
   BUFX2 U3087 ( .A(n3444), .Y(n2761));
   BUFX2 U3088 ( .A(n3316), .Y(n2762));
   BUFX2 U3089 ( .A(n3188), .Y(n2763));
   AND2X1 U3090 ( .A(w_mem_inst_N711),  .B(n3094), .Y(n3108));
   INVX1 U3091 ( .A(n3108), .Y(n2764));
   BUFX2 U3092 ( .A(n4945), .Y(n2765));
   BUFX2 U3093 ( .A(n5073), .Y(n2766));
   BUFX2 U3094 ( .A(n5189), .Y(n2767));
   BUFX2 U3095 ( .A(n5301), .Y(n2768));
   BUFX2 U3096 ( .A(n5353), .Y(n2769));
   BUFX2 U3097 ( .A(n5453), .Y(n2770));
   BUFX2 U3098 ( .A(n5583), .Y(n2771));
   BUFX2 U3099 ( .A(n5694), .Y(n2772));
   BUFX2 U3100 ( .A(n5720), .Y(n2773));
   BUFX2 U3101 ( .A(n4791), .Y(n2774));
   BUFX2 U3102 ( .A(n4829), .Y(n2775));
   INVX1 U3103 ( .A(n3103), .Y(n2776));
   BUFX2 U3104 ( .A(n3104), .Y(n2777));
   AND2X1 U3105 ( .A(n6067),  .B(t_ctr_reg[3]), .Y(n6089));
   INVX1 U3106 ( .A(n6089), .Y(n2778));
   BUFX2 U3107 ( .A(k_data[11]), .Y(n2779));
   AND2X2 U3108 ( .A(n6095),  .B(n6096), .Y(n6094));
   AND2X1 U3109 ( .A(n5771),  .B(n2893), .Y(n5912));
   INVX1 U3110 ( .A(n5912), .Y(n2780));
   AND2X1 U3111 ( .A(n5788),  .B(n4705), .Y(n5934));
   INVX1 U3112 ( .A(n5934), .Y(n2781));
   AND2X1 U3113 ( .A(t_ctr_reg[5]),  .B(n5998), .Y(n6000));
   INVX1 U3114 ( .A(n6000), .Y(n2782));
   AND2X1 U3115 ( .A(n6021),  .B(n4707), .Y(n5772));
   INVX1 U3116 ( .A(n5772), .Y(n2783));
   INVX1 U3117 ( .A(n5848), .Y(n2784));
   INVX1 U3118 ( .A(n5816), .Y(n2785));
   AND2X1 U3119 ( .A(N764),  .B(n3087), .Y(n5209));
   INVX1 U3120 ( .A(n5209), .Y(n2786));
   AND2X1 U3121 ( .A(N800),  .B(n3085), .Y(n5345));
   INVX1 U3122 ( .A(n5345), .Y(n2787));
   AND2X1 U3123 ( .A(N616),  .B(n3085), .Y(n5682));
   INVX1 U3124 ( .A(n5682), .Y(n2788));
   AND2X1 U3125 ( .A(N644),  .B(n3087), .Y(n5739));
   INVX1 U3126 ( .A(n5739), .Y(n2789));
   AND2X1 U3127 ( .A(N666),  .B(n3086), .Y(n4821));
   INVX1 U3128 ( .A(n4821), .Y(n2790));
   BUFX2 U3129 ( .A(n4124), .Y(n2791));
   BUFX2 U3130 ( .A(n3932), .Y(n2792));
   BUFX2 U3131 ( .A(n3740), .Y(n2793));
   BUFX2 U3132 ( .A(n3292), .Y(n2794));
   BUFX2 U3133 ( .A(n3164), .Y(n2795));
   BUFX2 U3134 ( .A(n3476), .Y(n2796));
   BUFX2 U3135 ( .A(n3794), .Y(n2797));
   BUFX2 U3136 ( .A(n3344), .Y(n2798));
   BUFX2 U3137 ( .A(n3216), .Y(n2799));
   BUFX2 U3138 ( .A(n3980), .Y(n2800));
   BUFX2 U3139 ( .A(n3596), .Y(n2801));
   BUFX2 U3140 ( .A(n3404), .Y(n2802));
   BUFX2 U3141 ( .A(n4042), .Y(n2803));
   BUFX2 U3142 ( .A(n3848), .Y(n2804));
   BUFX2 U3143 ( .A(n3656), .Y(n2805));
   BUFX2 U3144 ( .A(n3528), .Y(n2806));
   BUFX2 U3145 ( .A(n3142), .Y(n2807));
   BUFX2 U3146 ( .A(n4100), .Y(n2808));
   BUFX2 U3147 ( .A(n3908), .Y(n2809));
   BUFX2 U3148 ( .A(n3716), .Y(n2810));
   BUFX2 U3149 ( .A(n3450), .Y(n2811));
   BUFX2 U3150 ( .A(n4086), .Y(n2812));
   BUFX2 U3151 ( .A(n3958), .Y(n2813));
   BUFX2 U3152 ( .A(n3830), .Y(n2814));
   BUFX2 U3153 ( .A(n3702), .Y(n2815));
   BUFX2 U3154 ( .A(n3574), .Y(n2816));
   BUFX2 U3155 ( .A(n3446), .Y(n2817));
   BUFX2 U3156 ( .A(n3318), .Y(n2818));
   BUFX2 U3157 ( .A(n3190), .Y(n2819));
   BUFX2 U3158 ( .A(n4020), .Y(n2820));
   BUFX2 U3159 ( .A(n3892), .Y(n2821));
   BUFX2 U3160 ( .A(n3764), .Y(n2822));
   BUFX2 U3161 ( .A(n3636), .Y(n2823));
   BUFX2 U3162 ( .A(n3508), .Y(n2824));
   BUFX2 U3163 ( .A(n3380), .Y(n2825));
   BUFX2 U3164 ( .A(n3252), .Y(n2826));
   BUFX2 U3165 ( .A(n3124), .Y(n2827));
   BUFX2 U3166 ( .A(n4947), .Y(n2828));
   BUFX2 U3167 ( .A(n5085), .Y(n2829));
   BUFX2 U3168 ( .A(n5193), .Y(n2830));
   BUFX2 U3169 ( .A(n5309), .Y(n2831));
   BUFX2 U3170 ( .A(n5423), .Y(n2832));
   BUFX2 U3171 ( .A(n5459), .Y(n2833));
   BUFX2 U3172 ( .A(n5585), .Y(n2834));
   BUFX2 U3173 ( .A(n5690), .Y(n2835));
   BUFX2 U3174 ( .A(n5730), .Y(n2836));
   BUFX2 U3175 ( .A(n4797), .Y(n2837));
   BUFX2 U3176 ( .A(n4833), .Y(n2838));
   AND2X1 U3177 ( .A(N709),  .B(n3086), .Y(n4971));
   INVX1 U3178 ( .A(n4971), .Y(n2839));
   AND2X1 U3179 ( .A(n3099),  .B(n3100), .Y(n3096));
   INVX1 U3180 ( .A(n3096), .Y(n2840));
   AND2X1 U3181 ( .A(w_mem_inst_add_1008_carry[5]),  .B(n3094), .Y(n3097));
   INVX1 U3182 ( .A(n3097), .Y(n2841));
   AND2X1 U3183 ( .A(n5831),  .B(n4703), .Y(n5843));
   INVX1 U3184 ( .A(n5843), .Y(n2842));
   AND2X1 U3185 ( .A(n5860),  .B(n4711), .Y(n5918));
   INVX1 U3186 ( .A(n5918), .Y(n2843));
   AND2X1 U3187 ( .A(t_ctr_reg[3]),  .B(t_ctr_reg[4]), .Y(n5885));
   INVX1 U3188 ( .A(n5885), .Y(n2844));
   AND2X1 U3189 ( .A(n5874),  .B(n5763), .Y(n6002));
   INVX1 U3190 ( .A(n6002), .Y(n2845));
   INVX1 U3191 ( .A(n5749), .Y(n2846));
   AND2X1 U3192 ( .A(n6118),  .B(n4705), .Y(n5771));
   INVX1 U3193 ( .A(n5771), .Y(n2847));
   INVX1 U3194 ( .A(n5793), .Y(n2848));
   AND2X1 U3195 ( .A(n4700),  .B(n4701), .Y(n5789));
   INVX1 U3196 ( .A(n5789), .Y(n2849));
   BUFX2 U3197 ( .A(n4122), .Y(n2850));
   BUFX2 U3198 ( .A(n3930), .Y(n2851));
   BUFX2 U3199 ( .A(n3738), .Y(n2852));
   BUFX2 U3200 ( .A(n3354), .Y(n2853));
   BUFX2 U3201 ( .A(n3474), .Y(n2854));
   BUFX2 U3202 ( .A(n3978), .Y(n2855));
   BUFX2 U3203 ( .A(n3594), .Y(n2856));
   BUFX2 U3204 ( .A(n3402), .Y(n2857));
   BUFX2 U3205 ( .A(n3210), .Y(n2858));
   BUFX2 U3206 ( .A(n4040), .Y(n2859));
   BUFX2 U3207 ( .A(n3784), .Y(n2860));
   BUFX2 U3208 ( .A(n3846), .Y(n2861));
   BUFX2 U3209 ( .A(n3654), .Y(n2862));
   BUFX2 U3210 ( .A(n3526), .Y(n2863));
   BUFX2 U3211 ( .A(n3270), .Y(n2864));
   BUFX2 U3212 ( .A(n3140), .Y(n2865));
   BUFX2 U3213 ( .A(n4098), .Y(n2866));
   BUFX2 U3214 ( .A(n3906), .Y(n2867));
   BUFX2 U3215 ( .A(n3714), .Y(n2868));
   BUFX2 U3216 ( .A(n3330), .Y(n2869));
   BUFX2 U3217 ( .A(n4018), .Y(n2870));
   BUFX2 U3218 ( .A(n3890), .Y(n2871));
   BUFX2 U3219 ( .A(n3762), .Y(n2872));
   BUFX2 U3220 ( .A(n3634), .Y(n2873));
   BUFX2 U3221 ( .A(n3506), .Y(n2874));
   BUFX2 U3222 ( .A(n3378), .Y(n2875));
   BUFX2 U3223 ( .A(n3250), .Y(n2876));
   BUFX2 U3224 ( .A(n3122), .Y(n2877));
   BUFX2 U3225 ( .A(n4080), .Y(n2878));
   BUFX2 U3226 ( .A(n3952), .Y(n2879));
   BUFX2 U3227 ( .A(n3824), .Y(n2880));
   BUFX2 U3228 ( .A(n3696), .Y(n2881));
   BUFX2 U3229 ( .A(n3568), .Y(n2882));
   BUFX2 U3230 ( .A(n3440), .Y(n2883));
   BUFX2 U3231 ( .A(n3312), .Y(n2884));
   BUFX2 U3232 ( .A(n3184), .Y(n2885));
   AND2X1 U3233 ( .A(w_mem_inst_N714),  .B(n3094), .Y(n3114));
   INVX1 U3234 ( .A(n3114), .Y(n2886));
   BUFX2 U3235 ( .A(n4696), .Y(n2887));
   AND2X1 U3236 ( .A(t_ctr_reg[4]),  .B(t_ctr_reg[2]), .Y(n5998));
   INVX1 U3237 ( .A(n5998), .Y(n2888));
   AND2X1 U3238 ( .A(n5885),  .B(t_ctr_reg[5]), .Y(n5831));
   INVX1 U3239 ( .A(n5831), .Y(n2889));
   AND2X1 U3240 ( .A(n5805),  .B(t_ctr_reg[3]), .Y(n5874));
   INVX1 U3241 ( .A(n5874), .Y(n2890));
   AND2X1 U3242 ( .A(t_ctr_reg[1]),  .B(n4700), .Y(n5917));
   INVX1 U3243 ( .A(n5917), .Y(n2891));
   AND2X1 U3244 ( .A(n6117),  .B(n4711), .Y(n5782));
   INVX1 U3245 ( .A(n5782), .Y(n2892));
   INVX1 U3246 ( .A(n5751), .Y(n2893));
   BUFX2 U3247 ( .A(n4445), .Y(n2894));
   AND2X1 U3248 ( .A(n4144),  .B(w_mem_inst_w_ctr_reg[3]), .Y(n4442));
   INVX1 U3249 ( .A(n4442), .Y(n2895));
   AND2X1 U3250 ( .A(N694),  .B(n3085), .Y(n4941));
   INVX1 U3251 ( .A(n4941), .Y(n2896));
   AND2X1 U3252 ( .A(N748),  .B(n3087), .Y(n5177));
   INVX1 U3253 ( .A(n5177), .Y(n2897));
   AND2X1 U3254 ( .A(N639),  .B(n3087), .Y(n5728));
   INVX1 U3255 ( .A(n5728), .Y(n2898));
   BUFX2 U3256 ( .A(n4120), .Y(n2899));
   BUFX2 U3257 ( .A(n3928), .Y(n2900));
   BUFX2 U3258 ( .A(n3736), .Y(n2901));
   BUFX2 U3259 ( .A(n3352), .Y(n2902));
   BUFX2 U3260 ( .A(n3792), .Y(n2903));
   BUFX2 U3261 ( .A(n3472), .Y(n2904));
   BUFX2 U3262 ( .A(n3976), .Y(n2905));
   BUFX2 U3263 ( .A(n3592), .Y(n2906));
   BUFX2 U3264 ( .A(n3400), .Y(n2907));
   BUFX2 U3265 ( .A(n3208), .Y(n2908));
   BUFX2 U3266 ( .A(n4038), .Y(n2909));
   BUFX2 U3267 ( .A(n3844), .Y(n2910));
   BUFX2 U3268 ( .A(n3652), .Y(n2911));
   BUFX2 U3269 ( .A(n3524), .Y(n2912));
   BUFX2 U3270 ( .A(n3268), .Y(n2913));
   BUFX2 U3271 ( .A(n3138), .Y(n2914));
   BUFX2 U3272 ( .A(n4096), .Y(n2915));
   BUFX2 U3273 ( .A(n3904), .Y(n2916));
   BUFX2 U3274 ( .A(n3712), .Y(n2917));
   BUFX2 U3275 ( .A(n3328), .Y(n2918));
   BUFX2 U3276 ( .A(n3448), .Y(n2919));
   BUFX2 U3277 ( .A(n4082), .Y(n2920));
   BUFX2 U3278 ( .A(n3954), .Y(n2921));
   BUFX2 U3279 ( .A(n3826), .Y(n2922));
   BUFX2 U3280 ( .A(n3698), .Y(n2923));
   BUFX2 U3281 ( .A(n3570), .Y(n2924));
   BUFX2 U3282 ( .A(n3442), .Y(n2925));
   BUFX2 U3283 ( .A(n3314), .Y(n2926));
   BUFX2 U3284 ( .A(n3186), .Y(n2927));
   BUFX2 U3285 ( .A(n4016), .Y(n2928));
   BUFX2 U3286 ( .A(n3888), .Y(n2929));
   BUFX2 U3287 ( .A(n3760), .Y(n2930));
   BUFX2 U3288 ( .A(n3632), .Y(n2931));
   BUFX2 U3289 ( .A(n3504), .Y(n2932));
   BUFX2 U3290 ( .A(n3376), .Y(n2933));
   BUFX2 U3291 ( .A(n3248), .Y(n2934));
   BUFX2 U3292 ( .A(n3119), .Y(n2935));
   BUFX2 U3293 ( .A(n5087), .Y(n2936));
   BUFX2 U3294 ( .A(n5195), .Y(n2937));
   BUFX2 U3295 ( .A(n5313), .Y(n2938));
   BUFX2 U3296 ( .A(n5347), .Y(n2939));
   BUFX2 U3297 ( .A(n5441), .Y(n2940));
   BUFX2 U3298 ( .A(n5591), .Y(n2941));
   BUFX2 U3299 ( .A(n5696), .Y(n2942));
   BUFX2 U3300 ( .A(n5736), .Y(n2943));
   BUFX2 U3301 ( .A(n4801), .Y(n2944));
   BUFX2 U3302 ( .A(n4839), .Y(n2945));
   AND2X1 U3303 ( .A(N773),  .B(n3086), .Y(n5227));
   INVX1 U3304 ( .A(n5227), .Y(n2946));
   AND2X1 U3305 ( .A(N805),  .B(n3086), .Y(n5355));
   INVX1 U3306 ( .A(n5355), .Y(n2947));
   AND2X1 U3307 ( .A(N581),  .B(n3087), .Y(n5483));
   INVX1 U3308 ( .A(n5483), .Y(n2948));
   AND2X1 U3309 ( .A(N645),  .B(n3086), .Y(n5741));
   INVX1 U3310 ( .A(n5741), .Y(n2949));
   AND2X1 U3311 ( .A(n2980),  .B(w_mem_inst_sha256_w_mem_ctrl_reg_0_), .Y(n3094));
   INVX1 U3312 ( .A(n3094), .Y(n2950));
   BUFX2 U3313 ( .A(n5737), .Y(n2951));
   AND2X1 U3314 ( .A(n6061),  .B(n5917), .Y(n6045));
   INVX1 U3315 ( .A(n6045), .Y(n2952));
   AND2X1 U3316 ( .A(n5859),  .B(t_ctr_reg[2]), .Y(n5814));
   INVX1 U3317 ( .A(n5814), .Y(n2953));
   AND2X1 U3318 ( .A(n6118),  .B(t_ctr_reg[3]), .Y(n5845));
   INVX1 U3319 ( .A(n5845), .Y(n2954));
   INVX1 U3320 ( .A(n5861), .Y(puf_7_wire_3));
   INVX1 U3321 ( .A(n5786), .Y(n2956));
   AND2X1 U3322 ( .A(n3098),  .B(n3113), .Y(n4144));
   INVX1 U3323 ( .A(n4144), .Y(n2957));
   BUFX2 U3324 ( .A(n4168), .Y(n2958));
   INVX1 U3325 ( .A(n1759), .Y(n3089));
   INVX1 U3326 ( .A(n1759), .Y(n3088));
   INVX1 U3327 ( .A(n3081), .Y(n3062));
   INVX1 U3328 ( .A(n3081), .Y(n3055));
   INVX1 U3329 ( .A(n3081), .Y(n3059));
   INVX1 U3330 ( .A(n3081), .Y(n3053));
   INVX1 U3331 ( .A(n3081), .Y(n3061));
   INVX1 U3332 ( .A(n3081), .Y(n3054));
   INVX1 U3333 ( .A(n3081), .Y(n3058));
   INVX1 U3334 ( .A(n3081), .Y(n3063));
   INVX1 U3335 ( .A(n3081), .Y(n3060));
   INVX1 U3336 ( .A(n3081), .Y(n3057));
   INVX1 U3337 ( .A(n3081), .Y(n3056));
   INVX1 U3338 ( .A(n3081), .Y(n3052));
   INVX1 U3339 ( .A(n3081), .Y(n3051));
   INVX1 U3340 ( .A(n3081), .Y(n3078));
   INVX1 U3341 ( .A(n3081), .Y(n3070));
   INVX1 U3342 ( .A(n3081), .Y(n3075));
   INVX1 U3343 ( .A(n3081), .Y(n3067));
   INVX1 U3344 ( .A(n3081), .Y(n3080));
   INVX1 U3345 ( .A(n3081), .Y(n3072));
   INVX1 U3346 ( .A(n3081), .Y(n3064));
   INVX1 U3347 ( .A(n3081), .Y(n3077));
   INVX1 U3348 ( .A(n3081), .Y(n3069));
   INVX1 U3349 ( .A(n3081), .Y(n3074));
   INVX1 U3350 ( .A(n3081), .Y(n3066));
   INVX1 U3351 ( .A(n3081), .Y(n3079));
   INVX1 U3352 ( .A(n3081), .Y(n3076));
   INVX1 U3353 ( .A(n3081), .Y(n3073));
   INVX1 U3354 ( .A(n3081), .Y(n3071));
   INVX1 U3355 ( .A(n3081), .Y(n3068));
   INVX1 U3356 ( .A(n3081), .Y(n3065));
   INVX1 U3357 ( .A(n3012), .Y(n3009));
   INVX1 U3358 ( .A(n3012), .Y(n3001));
   INVX1 U3359 ( .A(n3012), .Y(n2993));
   INVX1 U3360 ( .A(n3012), .Y(n3006));
   INVX1 U3361 ( .A(n3012), .Y(n2998));
   INVX1 U3362 ( .A(n3012), .Y(n2990));
   INVX1 U3363 ( .A(n3012), .Y(n3011));
   INVX1 U3364 ( .A(n3012), .Y(n3003));
   INVX1 U3365 ( .A(n3012), .Y(n2995));
   INVX1 U3366 ( .A(n3012), .Y(n2987));
   INVX1 U3367 ( .A(n3012), .Y(n3008));
   INVX1 U3368 ( .A(n3012), .Y(n3000));
   INVX1 U3369 ( .A(n3012), .Y(n2992));
   INVX1 U3370 ( .A(n3012), .Y(n3005));
   INVX1 U3371 ( .A(n3012), .Y(n2997));
   INVX1 U3372 ( .A(n3012), .Y(n2989));
   INVX1 U3373 ( .A(n3012), .Y(n3010));
   INVX1 U3374 ( .A(n3012), .Y(n3007));
   INVX1 U3375 ( .A(n3012), .Y(n3004));
   INVX1 U3376 ( .A(n3012), .Y(n3002));
   INVX1 U3377 ( .A(n3012), .Y(n2999));
   INVX1 U3378 ( .A(n3012), .Y(n2996));
   INVX1 U3379 ( .A(n3012), .Y(n2994));
   INVX1 U3380 ( .A(n3012), .Y(n2991));
   INVX1 U3381 ( .A(n3012), .Y(n2988));
   INVX1 U3382 ( .A(n3012), .Y(n2986));
   INVX1 U3383 ( .A(n3012), .Y(n2985));
   INVX1 U3384 ( .A(n3012), .Y(n2982));
   INVX1 U3385 ( .A(n3012), .Y(n2984));
   INVX1 U3386 ( .A(n3012), .Y(n2981));
   INVX1 U3387 ( .A(n3012), .Y(n2983));
   INVX1 U3388 ( .A(n2102), .Y(n2977));
   INVX1 U3389 ( .A(n2102), .Y(n2979));
   INVX1 U3390 ( .A(n2102), .Y(n2978));
   INVX1 U3391 ( .A(n3049), .Y(n3016));
   INVX1 U3392 ( .A(n3049), .Y(n3015));
   INVX1 U3393 ( .A(n2102), .Y(n2980));
   INVX1 U3394 ( .A(n1852), .Y(n3027));
   INVX1 U3395 ( .A(n3049), .Y(n3032));
   INVX1 U3396 ( .A(n1852), .Y(n3039));
   INVX1 U3397 ( .A(n1852), .Y(n3017));
   INVX1 U3398 ( .A(n1852), .Y(n3022));
   INVX1 U3399 ( .A(n1852), .Y(n3038));
   INVX1 U3400 ( .A(n1852), .Y(n3025));
   INVX1 U3401 ( .A(n3049), .Y(n3030));
   INVX1 U3402 ( .A(n1852), .Y(n3042));
   INVX1 U3403 ( .A(n1852), .Y(n3035));
   INVX1 U3404 ( .A(n3049), .Y(n3020));
   INVX1 U3405 ( .A(n3049), .Y(n3028));
   INVX1 U3406 ( .A(n1852), .Y(n3033));
   INVX1 U3407 ( .A(n1852), .Y(n3018));
   INVX1 U3408 ( .A(n1852), .Y(n3040));
   INVX1 U3409 ( .A(n1852), .Y(n3023));
   INVX1 U3410 ( .A(n1852), .Y(n3037));
   INVX1 U3411 ( .A(n3049), .Y(n3026));
   INVX1 U3412 ( .A(n1852), .Y(n3029));
   INVX1 U3413 ( .A(n1852), .Y(n3031));
   INVX1 U3414 ( .A(n1852), .Y(n3034));
   INVX1 U3415 ( .A(n3049), .Y(n3019));
   INVX1 U3416 ( .A(n1852), .Y(n3021));
   INVX1 U3417 ( .A(n3049), .Y(n3024));
   INVX1 U3418 ( .A(n1852), .Y(n3041));
   INVX1 U3419 ( .A(n1852), .Y(n3036));
   INVX1 U3420 ( .A(n2887), .Y(n3085));
   INVX1 U3421 ( .A(n2887), .Y(n3086));
   INVX1 U3422 ( .A(n1852), .Y(n3045));
   INVX1 U3423 ( .A(n1852), .Y(n3043));
   INVX1 U3424 ( .A(n1852), .Y(n3044));
   INVX1 U3425 ( .A(n3049), .Y(n3046));
   INVX1 U3426 ( .A(n2887), .Y(n3087));
   INVX1 U3427 ( .A(n1852), .Y(n3047));
   INVX1 U3428 ( .A(n3049), .Y(n3048));
   INVX1 U3429 ( .A(n3092), .Y(n3093));
   INVX1 U3430 ( .A(n3120), .Y(n3081));
   INVX1 U3431 ( .A(n3084), .Y(n3083));
   INVX1 U3432 ( .A(n3084), .Y(n3082));
   INVX1 U3433 ( .A(n3049), .Y(n3013));
   INVX1 U3434 ( .A(n3049), .Y(n3014));
   INVX1 U3435 ( .A(n3050), .Y(n3049));
   AND2X1 U3436 ( .A(N902),  .B(N934), .Y(n2959));
   INVX1 U3437 ( .A(n4713), .Y(n3084));
   INVX1 U3438 ( .A(n2976), .Y(n3091));
   INVX1 U3439 ( .A(n2976), .Y(n3090));
   AND2X1 U3440 ( .A(t2[0]),  .B(N1029), .Y(n2960));
   AND2X1 U3441 ( .A(N870),  .B(k_data[0]), .Y(n2961));
   AND2X1 U3442 ( .A(w_mem_inst_N640),  .B(w_mem_inst_N672), .Y(n2962));
   INVX1 U3443 ( .A(n4783), .Y(n3092));
   INVX1 U3444 ( .A(n3117), .Y(n3012));
   AND2X1 U3445 ( .A(t1[0]),  .B(N997), .Y(n2963));
   AND2X1 U3446 ( .A(w_mem_inst_w_mem[192]),  .B(w_mem_inst_N639), .Y(n2964));
   AND2X1 U3447 ( .A(w_mem_inst_w_mem[480]),  .B(w_mem_inst_N607), .Y(n2965));
   AND2X1 U3448 ( .A(N837),  .B(h_reg[0]), .Y(n2966));
   AND2X1 U3449 ( .A(t1[0]),  .B(d_reg[0]), .Y(n2967));
   AND2X1 U3450 ( .A(b_reg[0]),  .B(digest[192]), .Y(n2968));
   AND2X1 U3451 ( .A(h_reg[0]),  .B(digest[0]), .Y(n2969));
   AND2X1 U3452 ( .A(f_reg[0]),  .B(digest[64]), .Y(n2970));
   AND2X1 U3453 ( .A(d_reg[0]),  .B(digest[128]), .Y(n2971));
   AND2X1 U3454 ( .A(c_reg[0]),  .B(digest[160]), .Y(n2972));
   AND2X1 U3455 ( .A(a_reg[0]),  .B(digest[224]), .Y(n2973));
   AND2X1 U3456 ( .A(g_reg[0]),  .B(digest[32]), .Y(n2974));
   AND2X1 U3457 ( .A(e_reg[0]),  .B(digest[96]), .Y(n2975));
   AND2X1 U3458 ( .A(init),  .B(n3046), .Y(n2976));
   INVX1 U3459 ( .A(n1852), .Y(n3050));
   XOR2X1 U3460 ( .A(w_mem_inst_w_mem[192]),  .B(w_mem_inst_N639), .Y(w_mem_inst_N640));
   XOR2X1 U3461 ( .A(w_mem_inst_w_mem[480]),  .B(w_mem_inst_N607), .Y(w_mem_inst_N672));
   XOR2X1 U3462 ( .A(w_mem_inst_N672),  .B(w_mem_inst_N640), .Y(w_mem_inst_w_new[0]));
   XOR2X1 U3463 ( .A(t1[0]),  .B(d_reg[0]), .Y(N1579));
   XOR2X1 U3464 ( .A(t2[0]),  .B(N1029), .Y(N1547));
   XOR2X1 U3465 ( .A(N997),  .B(t1[0]), .Y(t2[0]));
   XOR2X1 U3466 ( .A(N934),  .B(N902), .Y(t1[0]));
   XOR2X1 U3467 ( .A(N870),  .B(k_data[0]), .Y(N934));
   XOR2X1 U3468 ( .A(n1849),  .B(N869), .Y(N902));
   XOR2X1 U3469 ( .A(N837),  .B(h_reg[0]), .Y(N870));
   XOR2X1 U3470 ( .A(h_reg[0]),  .B(digest[0]), .Y(N774));
   XOR2X1 U3471 ( .A(g_reg[0]),  .B(digest[32]), .Y(N742));
   XOR2X1 U3472 ( .A(f_reg[0]),  .B(digest[64]), .Y(N710));
   XOR2X1 U3473 ( .A(e_reg[0]),  .B(digest[96]), .Y(N678));
   XOR2X1 U3474 ( .A(d_reg[0]),  .B(digest[128]), .Y(N646));
   XOR2X1 U3475 ( .A(c_reg[0]),  .B(digest[160]), .Y(N614));
   XOR2X1 U3476 ( .A(b_reg[0]),  .B(digest[192]), .Y(N582));
   XOR2X1 U3477 ( .A(a_reg[0]),  .B(digest[224]), .Y(N550));
   MUX2X1 U3478 ( .A(n3095),  .B(n2950),  .S(w_mem_inst_w_ctr_reg[0]), .Y(w_mem_inst_n2142));
   MUX2X1 U3479 ( .A(n2841),  .B(n2840),  .S(n3098), .Y(w_mem_inst_n2141));
   OAI21X1 U3480 ( .A(w_mem_inst_add_1008_carry[5]),  .B(n3101),  .C(n3102), .Y(n3099));
   MUX2X1 U3481 ( .A(n1852),  .B(n2776),  .S(n3101), .Y(w_mem_inst_n2140));
   NAND3X1 U3482 ( .A(w_mem_inst_w_ctr_reg[4]),  .B(w_mem_inst_w_ctr_reg[3]),  .C(n3105), .Y(n3104));
   AND2X1 U3483 ( .A(w_mem_inst_w_ctr_reg[5]),  .B(n3106), .Y(n3105));
   OAI21X1 U3484 ( .A(n3095),  .B(n3107),  .C(n2764), .Y(w_mem_inst_n2139));
   OAI21X1 U3485 ( .A(n3095),  .B(n3109),  .C(n2701), .Y(w_mem_inst_n2138));
   OAI21X1 U3486 ( .A(n3095),  .B(n3111),  .C(n2638), .Y(w_mem_inst_n2137));
   OAI21X1 U3487 ( .A(n3095),  .B(n3113),  .C(n2886), .Y(w_mem_inst_n2136));
   OR2X1 U3488 ( .A(n3102),  .B(rst), .Y(n3095));
   MUX2X1 U3489 ( .A(n3116),  .B(n1958),  .S(n3101), .Y(n3102));
   INVX1 U3490 ( .A(w_mem_inst_sha256_w_mem_ctrl_reg_0_), .Y(n3101));
   OAI21X1 U3491 ( .A(n3007),  .B(n3118),  .C(n2935), .Y(w_mem_inst_n2135));
   AOI22X1 U3492 ( .A(block[0]),  .B(n3039),  .C(w_mem_inst_w_new[0]),  .D(n3120), .Y(n3119));
   OAI21X1 U3493 ( .A(n2993),  .B(n3121),  .C(n2877), .Y(w_mem_inst_n2134));
   AOI22X1 U3494 ( .A(block[1]),  .B(n3013),  .C(w_mem_inst_w_new[1]),  .D(n3120), .Y(n3122));
   OAI21X1 U3495 ( .A(n2981),  .B(n3123),  .C(n2827), .Y(w_mem_inst_n2133));
   AOI22X1 U3496 ( .A(block[2]),  .B(n3030),  .C(w_mem_inst_w_new[2]),  .D(n3120), .Y(n3124));
   INVX1 U3497 ( .A(w_mem_inst_w_mem[2]), .Y(n3123));
   OAI21X1 U3498 ( .A(n2992),  .B(n3125),  .C(n2755), .Y(w_mem_inst_n2132));
   AOI22X1 U3499 ( .A(block[3]),  .B(n3024),  .C(w_mem_inst_w_new[3]),  .D(n3120), .Y(n3126));
   INVX1 U3500 ( .A(w_mem_inst_w_mem[3]), .Y(n3125));
   OAI21X1 U3501 ( .A(n3009),  .B(n3127),  .C(n2637), .Y(w_mem_inst_n2131));
   AOI22X1 U3502 ( .A(block[4]),  .B(n3024),  .C(w_mem_inst_w_new[4]),  .D(n3120), .Y(n3128));
   INVX1 U3503 ( .A(w_mem_inst_w_mem[4]), .Y(n3127));
   OAI21X1 U3504 ( .A(n2998),  .B(n3129),  .C(n2523), .Y(w_mem_inst_n2130));
   AOI22X1 U3505 ( .A(block[5]),  .B(n3024),  .C(w_mem_inst_w_new[5]),  .D(n3120), .Y(n3130));
   INVX1 U3506 ( .A(w_mem_inst_w_mem[5]), .Y(n3129));
   OAI21X1 U3507 ( .A(n2987),  .B(n3131),  .C(n2470), .Y(w_mem_inst_n2129));
   AOI22X1 U3508 ( .A(block[6]),  .B(n3024),  .C(w_mem_inst_w_new[6]),  .D(n3120), .Y(n3132));
   INVX1 U3509 ( .A(w_mem_inst_w_mem[6]), .Y(n3131));
   OAI21X1 U3510 ( .A(n2994),  .B(n3133),  .C(n2414), .Y(w_mem_inst_n2128));
   AOI22X1 U3511 ( .A(block[7]),  .B(n3024),  .C(w_mem_inst_w_new[7]),  .D(n3120), .Y(n3134));
   INVX1 U3512 ( .A(w_mem_inst_w_mem[7]), .Y(n3133));
   OAI21X1 U3513 ( .A(n3011),  .B(n3135),  .C(n2358), .Y(w_mem_inst_n2127));
   AOI22X1 U3514 ( .A(block[8]),  .B(n3024),  .C(w_mem_inst_w_new[8]),  .D(n3080), .Y(n3136));
   INVX1 U3515 ( .A(w_mem_inst_w_mem[8]), .Y(n3135));
   OAI21X1 U3516 ( .A(n3011),  .B(n3137),  .C(n2914), .Y(w_mem_inst_n2126));
   AOI22X1 U3517 ( .A(block[9]),  .B(n3025),  .C(w_mem_inst_w_new[9]),  .D(n3080), .Y(n3138));
   INVX1 U3518 ( .A(w_mem_inst_w_mem[9]), .Y(n3137));
   OAI21X1 U3519 ( .A(n3011),  .B(n3139),  .C(n2865), .Y(w_mem_inst_n2125));
   AOI22X1 U3520 ( .A(block[10]),  .B(n3025),  .C(w_mem_inst_w_new[10]),  .D(n3080), .Y(n3140));
   OAI21X1 U3521 ( .A(n3011),  .B(n3141),  .C(n2807), .Y(w_mem_inst_n2124));
   AOI22X1 U3522 ( .A(block[11]),  .B(n3025),  .C(w_mem_inst_w_new[11]),  .D(n3080), .Y(n3142));
   OAI21X1 U3523 ( .A(n3011),  .B(n3143),  .C(n2743), .Y(w_mem_inst_n2123));
   AOI22X1 U3524 ( .A(block[12]),  .B(n3025),  .C(w_mem_inst_w_new[12]),  .D(n3080), .Y(n3144));
   OAI21X1 U3525 ( .A(n3011),  .B(n3145),  .C(n2684), .Y(w_mem_inst_n2122));
   AOI22X1 U3526 ( .A(block[13]),  .B(n3025),  .C(w_mem_inst_w_new[13]),  .D(n3080), .Y(n3146));
   OAI21X1 U3527 ( .A(n3011),  .B(n3147),  .C(n2621), .Y(w_mem_inst_n2121));
   AOI22X1 U3528 ( .A(block[14]),  .B(n3025),  .C(w_mem_inst_w_new[14]),  .D(n3080), .Y(n3148));
   OAI21X1 U3529 ( .A(n3011),  .B(n3149),  .C(n2565), .Y(w_mem_inst_n2120));
   AOI22X1 U3530 ( .A(block[15]),  .B(n3025),  .C(w_mem_inst_w_new[15]),  .D(n3080), .Y(n3150));
   OAI21X1 U3531 ( .A(n3011),  .B(n3151),  .C(n2507), .Y(w_mem_inst_n2119));
   AOI22X1 U3532 ( .A(block[16]),  .B(n3025),  .C(w_mem_inst_w_new[16]),  .D(n3080), .Y(n3152));
   OAI21X1 U3533 ( .A(n3011),  .B(n3153),  .C(n2454), .Y(w_mem_inst_n2118));
   AOI22X1 U3534 ( .A(block[17]),  .B(n3025),  .C(w_mem_inst_w_new[17]),  .D(n3080), .Y(n3154));
   OAI21X1 U3535 ( .A(n3011),  .B(n3155),  .C(n2398), .Y(w_mem_inst_n2117));
   AOI22X1 U3536 ( .A(block[18]),  .B(n3025),  .C(w_mem_inst_w_new[18]),  .D(n3080), .Y(n3156));
   OAI21X1 U3537 ( .A(n3011),  .B(n3157),  .C(n2290), .Y(w_mem_inst_n2116));
   AOI22X1 U3538 ( .A(block[19]),  .B(n3025),  .C(w_mem_inst_w_new[19]),  .D(n3080), .Y(n3158));
   OAI21X1 U3539 ( .A(n3010),  .B(n3159),  .C(n2342), .Y(w_mem_inst_n2115));
   AOI22X1 U3540 ( .A(block[20]),  .B(n3025),  .C(w_mem_inst_w_new[20]),  .D(n3079), .Y(n3160));
   OAI21X1 U3541 ( .A(n3010),  .B(n3161),  .C(n2247), .Y(w_mem_inst_n2114));
   AOI22X1 U3542 ( .A(block[21]),  .B(n3025),  .C(w_mem_inst_w_new[21]),  .D(n3079), .Y(n3162));
   OAI21X1 U3543 ( .A(n3010),  .B(n3163),  .C(n2795), .Y(w_mem_inst_n2113));
   AOI22X1 U3544 ( .A(block[22]),  .B(n3026),  .C(w_mem_inst_w_new[22]),  .D(n3079), .Y(n3164));
   OAI21X1 U3545 ( .A(n3010),  .B(n3165),  .C(n2669), .Y(w_mem_inst_n2112));
   AOI22X1 U3546 ( .A(block[23]),  .B(n3026),  .C(w_mem_inst_w_new[23]),  .D(n3079), .Y(n3166));
   INVX1 U3547 ( .A(w_mem_inst_w_mem[23]), .Y(n3165));
   OAI21X1 U3548 ( .A(n3010),  .B(n3167),  .C(n2605), .Y(w_mem_inst_n2111));
   AOI22X1 U3549 ( .A(block[24]),  .B(n3026),  .C(w_mem_inst_w_new[24]),  .D(n3079), .Y(n3168));
   INVX1 U3550 ( .A(w_mem_inst_w_mem[24]), .Y(n3167));
   OAI21X1 U3551 ( .A(n3010),  .B(n3169),  .C(n2550), .Y(w_mem_inst_n2110));
   AOI22X1 U3552 ( .A(block[25]),  .B(n3026),  .C(w_mem_inst_w_new[25]),  .D(n3079), .Y(n3170));
   INVX1 U3553 ( .A(w_mem_inst_w_mem[25]), .Y(n3169));
   OAI21X1 U3554 ( .A(n3010),  .B(n3171),  .C(n2491), .Y(w_mem_inst_n2109));
   AOI22X1 U3555 ( .A(block[26]),  .B(n3026),  .C(w_mem_inst_w_new[26]),  .D(n3079), .Y(n3172));
   INVX1 U3556 ( .A(w_mem_inst_w_mem[26]), .Y(n3171));
   OAI21X1 U3557 ( .A(n3010),  .B(n3173),  .C(n2438), .Y(w_mem_inst_n2108));
   AOI22X1 U3558 ( .A(block[27]),  .B(n3026),  .C(w_mem_inst_w_new[27]),  .D(n3079), .Y(n3174));
   INVX1 U3559 ( .A(w_mem_inst_w_mem[27]), .Y(n3173));
   OAI21X1 U3560 ( .A(n3010),  .B(n3175),  .C(n2382), .Y(w_mem_inst_n2107));
   AOI22X1 U3561 ( .A(block[28]),  .B(n3026),  .C(w_mem_inst_w_new[28]),  .D(n3079), .Y(n3176));
   INVX1 U3562 ( .A(w_mem_inst_w_mem[28]), .Y(n3175));
   OAI21X1 U3563 ( .A(n3010),  .B(n3177),  .C(n2275), .Y(w_mem_inst_n2106));
   AOI22X1 U3564 ( .A(block[29]),  .B(n3026),  .C(w_mem_inst_w_new[29]),  .D(n3079), .Y(n3178));
   INVX1 U3565 ( .A(w_mem_inst_w_mem[29]), .Y(n3177));
   OAI21X1 U3566 ( .A(n3010),  .B(n3179),  .C(n2202), .Y(w_mem_inst_n2105));
   AOI22X1 U3567 ( .A(block[30]),  .B(n3026),  .C(w_mem_inst_w_new[30]),  .D(n3079), .Y(n3180));
   INVX1 U3568 ( .A(w_mem_inst_w_mem[30]), .Y(n3179));
   OAI21X1 U3569 ( .A(n3010),  .B(n3181),  .C(n2179), .Y(w_mem_inst_n2104));
   AOI22X1 U3570 ( .A(block[31]),  .B(n3026),  .C(w_mem_inst_w_new[31]),  .D(n3079), .Y(n3182));
   INVX1 U3571 ( .A(w_mem_inst_w_mem[31]), .Y(n3181));
   OAI21X1 U3572 ( .A(n3009),  .B(n3183),  .C(n2885), .Y(w_mem_inst_n2103));
   AOI22X1 U3573 ( .A(block[32]),  .B(n3026),  .C(w_mem_inst_w_mem[0]),  .D(n3078), .Y(n3184));
   OAI21X1 U3574 ( .A(n3009),  .B(n3185),  .C(n2927), .Y(w_mem_inst_n2102));
   AOI22X1 U3575 ( .A(block[33]),  .B(n3026),  .C(w_mem_inst_w_mem[1]),  .D(n3078), .Y(n3186));
   OAI21X1 U3576 ( .A(n3009),  .B(n3187),  .C(n2763), .Y(w_mem_inst_n2101));
   AOI22X1 U3577 ( .A(block[34]),  .B(n3026),  .C(w_mem_inst_w_mem[2]),  .D(n3078), .Y(n3188));
   OAI21X1 U3578 ( .A(n3009),  .B(n3189),  .C(n2819), .Y(w_mem_inst_n2100));
   AOI22X1 U3579 ( .A(block[35]),  .B(n3027),  .C(w_mem_inst_w_mem[3]),  .D(n3078), .Y(n3190));
   OAI21X1 U3580 ( .A(n3009),  .B(n3191),  .C(n2699), .Y(w_mem_inst_n2099));
   AOI22X1 U3581 ( .A(block[36]),  .B(n3027),  .C(w_mem_inst_w_mem[4]),  .D(n3078), .Y(n3192));
   OAI21X1 U3582 ( .A(n3009),  .B(n3193),  .C(n2630), .Y(w_mem_inst_n2098));
   AOI22X1 U3583 ( .A(block[37]),  .B(n3027),  .C(w_mem_inst_w_mem[5]),  .D(n3078), .Y(n3194));
   OAI21X1 U3584 ( .A(n3009),  .B(n3195),  .C(n2580), .Y(w_mem_inst_n2097));
   AOI22X1 U3585 ( .A(block[38]),  .B(n3027),  .C(w_mem_inst_w_mem[6]),  .D(n3078), .Y(n3196));
   OAI21X1 U3586 ( .A(n3009),  .B(n3197),  .C(n2516), .Y(w_mem_inst_n2096));
   AOI22X1 U3587 ( .A(block[39]),  .B(n3027),  .C(w_mem_inst_w_mem[7]),  .D(n3078), .Y(n3198));
   OAI21X1 U3588 ( .A(n3009),  .B(n3199),  .C(n2468), .Y(w_mem_inst_n2095));
   AOI22X1 U3589 ( .A(block[40]),  .B(n3027),  .C(w_mem_inst_w_mem[8]),  .D(n3078), .Y(n3200));
   OAI21X1 U3590 ( .A(n3009),  .B(n3201),  .C(n2410), .Y(w_mem_inst_n2094));
   AOI22X1 U3591 ( .A(block[41]),  .B(n3027),  .C(w_mem_inst_w_mem[9]),  .D(n3078), .Y(n3202));
   OAI21X1 U3592 ( .A(n3009),  .B(n3203),  .C(n2356), .Y(w_mem_inst_n2093));
   AOI22X1 U3593 ( .A(block[42]),  .B(n3027),  .C(w_mem_inst_w_mem[10]),  .D(n3078), .Y(n3204));
   OAI21X1 U3594 ( .A(n3009),  .B(n3205),  .C(n2303), .Y(w_mem_inst_n2092));
   AOI22X1 U3595 ( .A(block[43]),  .B(n3027),  .C(w_mem_inst_w_mem[11]),  .D(n3078), .Y(n3206));
   OAI21X1 U3596 ( .A(n3008),  .B(n3207),  .C(n2908), .Y(w_mem_inst_n2091));
   AOI22X1 U3597 ( .A(block[44]),  .B(n3027),  .C(w_mem_inst_w_mem[12]),  .D(n3077), .Y(n3208));
   OAI21X1 U3598 ( .A(n3008),  .B(n3209),  .C(n2858), .Y(w_mem_inst_n2090));
   AOI22X1 U3599 ( .A(block[45]),  .B(n3027),  .C(w_mem_inst_w_mem[13]),  .D(n3077), .Y(n3210));
   OAI21X1 U3600 ( .A(n3008),  .B(n3211),  .C(n2739), .Y(w_mem_inst_n2089));
   AOI22X1 U3601 ( .A(block[46]),  .B(n3027),  .C(w_mem_inst_w_mem[14]),  .D(n3077), .Y(n3212));
   OAI21X1 U3602 ( .A(n3008),  .B(n3213),  .C(n2255), .Y(w_mem_inst_n2088));
   AOI22X1 U3603 ( .A(block[47]),  .B(n3027),  .C(w_mem_inst_w_mem[15]),  .D(n3077), .Y(n3214));
   OAI21X1 U3604 ( .A(n3008),  .B(n3215),  .C(n2799), .Y(w_mem_inst_n2087));
   AOI22X1 U3605 ( .A(block[48]),  .B(n3028),  .C(w_mem_inst_w_mem[16]),  .D(n3077), .Y(n3216));
   OAI21X1 U3606 ( .A(n3008),  .B(n3217),  .C(n2676), .Y(w_mem_inst_n2086));
   AOI22X1 U3607 ( .A(block[49]),  .B(n3028),  .C(w_mem_inst_w_mem[17]),  .D(n3077), .Y(n3218));
   OAI21X1 U3608 ( .A(n3008),  .B(n3219),  .C(n2614), .Y(w_mem_inst_n2085));
   AOI22X1 U3609 ( .A(block[50]),  .B(n3028),  .C(w_mem_inst_w_mem[18]),  .D(n3077), .Y(n3220));
   OAI21X1 U3610 ( .A(n3008),  .B(n3221),  .C(n2557), .Y(w_mem_inst_n2084));
   AOI22X1 U3611 ( .A(block[51]),  .B(n3028),  .C(w_mem_inst_w_mem[19]),  .D(n3077), .Y(n3222));
   OAI21X1 U3612 ( .A(n3008),  .B(n3223),  .C(n2500), .Y(w_mem_inst_n2083));
   AOI22X1 U3613 ( .A(block[52]),  .B(n3028),  .C(w_mem_inst_w_mem[20]),  .D(n3077), .Y(n3224));
   OAI21X1 U3614 ( .A(n3008),  .B(n3225),  .C(n2447), .Y(w_mem_inst_n2082));
   AOI22X1 U3615 ( .A(block[53]),  .B(n3028),  .C(w_mem_inst_w_mem[21]),  .D(n3077), .Y(n3226));
   OAI21X1 U3616 ( .A(n3008),  .B(n3227),  .C(n2392), .Y(w_mem_inst_n2081));
   AOI22X1 U3617 ( .A(block[54]),  .B(n3028),  .C(w_mem_inst_w_mem[22]),  .D(n3077), .Y(n3228));
   OAI21X1 U3618 ( .A(n3008),  .B(n3229),  .C(n2340), .Y(w_mem_inst_n2080));
   AOI22X1 U3619 ( .A(block[55]),  .B(n3028),  .C(w_mem_inst_w_mem[23]),  .D(n3077), .Y(n3230));
   OAI21X1 U3620 ( .A(n3007),  .B(n3231),  .C(n2285), .Y(w_mem_inst_n2079));
   AOI22X1 U3621 ( .A(block[56]),  .B(n3028),  .C(w_mem_inst_w_mem[24]),  .D(n3076), .Y(n3232));
   OAI21X1 U3622 ( .A(n3007),  .B(n3233),  .C(n2242), .Y(w_mem_inst_n2078));
   AOI22X1 U3623 ( .A(block[57]),  .B(n3028),  .C(w_mem_inst_w_mem[25]),  .D(n3076), .Y(n3234));
   OAI21X1 U3624 ( .A(n3007),  .B(n3235),  .C(n2209), .Y(w_mem_inst_n2077));
   AOI22X1 U3625 ( .A(block[58]),  .B(n3028),  .C(w_mem_inst_w_mem[26]),  .D(n3076), .Y(n3236));
   OAI21X1 U3626 ( .A(n3007),  .B(n3237),  .C(n2186), .Y(w_mem_inst_n2076));
   AOI22X1 U3627 ( .A(block[59]),  .B(n3028),  .C(w_mem_inst_w_mem[27]),  .D(n3076), .Y(n3238));
   OAI21X1 U3628 ( .A(n3007),  .B(n3239),  .C(n2164), .Y(w_mem_inst_n2075));
   AOI22X1 U3629 ( .A(block[60]),  .B(n3028),  .C(w_mem_inst_w_mem[28]),  .D(n3076), .Y(n3240));
   OAI21X1 U3630 ( .A(n3007),  .B(n3241),  .C(n2326), .Y(w_mem_inst_n2074));
   AOI22X1 U3631 ( .A(block[61]),  .B(n3029),  .C(w_mem_inst_w_mem[29]),  .D(n3076), .Y(n3242));
   OAI21X1 U3632 ( .A(n3007),  .B(n3243),  .C(n2149), .Y(w_mem_inst_n2073));
   AOI22X1 U3633 ( .A(block[62]),  .B(n3029),  .C(w_mem_inst_w_mem[30]),  .D(n3076), .Y(n3244));
   OAI21X1 U3634 ( .A(n3007),  .B(n3245),  .C(n2137), .Y(w_mem_inst_n2072));
   AOI22X1 U3635 ( .A(block[63]),  .B(n3029),  .C(w_mem_inst_w_mem[31]),  .D(n3076), .Y(n3246));
   OAI21X1 U3636 ( .A(n3007),  .B(n3247),  .C(n2934), .Y(w_mem_inst_n2071));
   AOI22X1 U3637 ( .A(block[64]),  .B(n3029),  .C(w_mem_inst_w_mem[32]),  .D(n3076), .Y(n3248));
   INVX1 U3638 ( .A(w_mem_inst_w_mem[64]), .Y(n3247));
   OAI21X1 U3639 ( .A(n3007),  .B(n3249),  .C(n2876), .Y(w_mem_inst_n2070));
   AOI22X1 U3640 ( .A(block[65]),  .B(n3029),  .C(w_mem_inst_w_mem[33]),  .D(n3076), .Y(n3250));
   INVX1 U3641 ( .A(w_mem_inst_w_mem[65]), .Y(n3249));
   OAI21X1 U3642 ( .A(n3007),  .B(n3251),  .C(n2826), .Y(w_mem_inst_n2069));
   AOI22X1 U3643 ( .A(block[66]),  .B(n3029),  .C(w_mem_inst_w_mem[34]),  .D(n3076), .Y(n3252));
   INVX1 U3644 ( .A(w_mem_inst_w_mem[66]), .Y(n3251));
   OAI21X1 U3645 ( .A(n3007),  .B(n3253),  .C(n2754), .Y(w_mem_inst_n2068));
   AOI22X1 U3646 ( .A(block[67]),  .B(n3029),  .C(w_mem_inst_w_mem[35]),  .D(n3076), .Y(n3254));
   INVX1 U3647 ( .A(w_mem_inst_w_mem[67]), .Y(n3253));
   OAI21X1 U3648 ( .A(n3006),  .B(n3255),  .C(n2636), .Y(w_mem_inst_n2067));
   AOI22X1 U3649 ( .A(block[68]),  .B(n3029),  .C(w_mem_inst_w_mem[36]),  .D(n3075), .Y(n3256));
   INVX1 U3650 ( .A(w_mem_inst_w_mem[68]), .Y(n3255));
   OAI21X1 U3651 ( .A(n3006),  .B(n3257),  .C(n2692), .Y(w_mem_inst_n2066));
   AOI22X1 U3652 ( .A(block[69]),  .B(n3029),  .C(w_mem_inst_w_mem[37]),  .D(n3075), .Y(n3258));
   INVX1 U3653 ( .A(w_mem_inst_w_mem[69]), .Y(n3257));
   OAI21X1 U3654 ( .A(n3006),  .B(n3259),  .C(n2522), .Y(w_mem_inst_n2065));
   AOI22X1 U3655 ( .A(block[70]),  .B(n3029),  .C(w_mem_inst_w_mem[38]),  .D(n3075), .Y(n3260));
   INVX1 U3656 ( .A(w_mem_inst_w_mem[70]), .Y(n3259));
   OAI21X1 U3657 ( .A(n3006),  .B(n3261),  .C(n2573), .Y(w_mem_inst_n2064));
   AOI22X1 U3658 ( .A(block[71]),  .B(n3029),  .C(w_mem_inst_w_mem[39]),  .D(n3075), .Y(n3262));
   INVX1 U3659 ( .A(w_mem_inst_w_mem[71]), .Y(n3261));
   OAI21X1 U3660 ( .A(n3006),  .B(n3263),  .C(n2413), .Y(w_mem_inst_n2063));
   AOI22X1 U3661 ( .A(block[72]),  .B(n3029),  .C(w_mem_inst_w_mem[40]),  .D(n3075), .Y(n3264));
   INVX1 U3662 ( .A(w_mem_inst_w_mem[72]), .Y(n3263));
   OAI21X1 U3663 ( .A(n3006),  .B(n3265),  .C(n2462), .Y(w_mem_inst_n2062));
   AOI22X1 U3664 ( .A(block[73]),  .B(n3029),  .C(w_mem_inst_w_mem[41]),  .D(n3075), .Y(n3266));
   INVX1 U3665 ( .A(w_mem_inst_w_mem[73]), .Y(n3265));
   OAI21X1 U3666 ( .A(n3006),  .B(n3267),  .C(n2913), .Y(w_mem_inst_n2061));
   AOI22X1 U3667 ( .A(block[74]),  .B(n3030),  .C(w_mem_inst_w_mem[42]),  .D(n3075), .Y(n3268));
   INVX1 U3668 ( .A(w_mem_inst_w_mem[74]), .Y(n3267));
   OAI21X1 U3669 ( .A(n3006),  .B(n3269),  .C(n2864), .Y(w_mem_inst_n2060));
   AOI22X1 U3670 ( .A(block[75]),  .B(n3030),  .C(w_mem_inst_w_mem[43]),  .D(n3075), .Y(n3270));
   INVX1 U3671 ( .A(w_mem_inst_w_mem[75]), .Y(n3269));
   OAI21X1 U3672 ( .A(n3006),  .B(n3271),  .C(n2742), .Y(w_mem_inst_n2059));
   AOI22X1 U3673 ( .A(block[76]),  .B(n3030),  .C(w_mem_inst_w_mem[44]),  .D(n3075), .Y(n3272));
   INVX1 U3674 ( .A(w_mem_inst_w_mem[76]), .Y(n3271));
   OAI21X1 U3675 ( .A(n3006),  .B(n3273),  .C(n2351), .Y(w_mem_inst_n2058));
   AOI22X1 U3676 ( .A(block[77]),  .B(n3030),  .C(w_mem_inst_w_mem[45]),  .D(n3075), .Y(n3274));
   INVX1 U3677 ( .A(w_mem_inst_w_mem[77]), .Y(n3273));
   OAI21X1 U3678 ( .A(n3006),  .B(n3275),  .C(n2297), .Y(w_mem_inst_n2057));
   AOI22X1 U3679 ( .A(block[78]),  .B(n3030),  .C(w_mem_inst_w_mem[46]),  .D(n3075), .Y(n3276));
   INVX1 U3680 ( .A(w_mem_inst_w_mem[78]), .Y(n3275));
   OAI21X1 U3681 ( .A(n3006),  .B(n3277),  .C(n2214), .Y(w_mem_inst_n2056));
   AOI22X1 U3682 ( .A(block[79]),  .B(n3030),  .C(w_mem_inst_w_mem[47]),  .D(n3075), .Y(n3278));
   INVX1 U3683 ( .A(w_mem_inst_w_mem[79]), .Y(n3277));
   OAI21X1 U3684 ( .A(n3005),  .B(n3279),  .C(n2681), .Y(w_mem_inst_n2055));
   AOI22X1 U3685 ( .A(block[80]),  .B(n3030),  .C(w_mem_inst_w_mem[48]),  .D(n3074), .Y(n3280));
   INVX1 U3686 ( .A(w_mem_inst_w_mem[80]), .Y(n3279));
   OAI21X1 U3687 ( .A(n3005),  .B(n3281),  .C(n2619), .Y(w_mem_inst_n2054));
   AOI22X1 U3688 ( .A(block[81]),  .B(n3030),  .C(w_mem_inst_w_mem[49]),  .D(n3074), .Y(n3282));
   INVX1 U3689 ( .A(w_mem_inst_w_mem[81]), .Y(n3281));
   OAI21X1 U3690 ( .A(n3005),  .B(n3283),  .C(n2562), .Y(w_mem_inst_n2053));
   AOI22X1 U3691 ( .A(block[82]),  .B(n3030),  .C(w_mem_inst_w_mem[50]),  .D(n3074), .Y(n3284));
   INVX1 U3692 ( .A(w_mem_inst_w_mem[82]), .Y(n3283));
   OAI21X1 U3693 ( .A(n3005),  .B(n3285),  .C(n2505), .Y(w_mem_inst_n2052));
   AOI22X1 U3694 ( .A(block[83]),  .B(n3030),  .C(w_mem_inst_w_mem[51]),  .D(n3074), .Y(n3286));
   INVX1 U3695 ( .A(w_mem_inst_w_mem[83]), .Y(n3285));
   OAI21X1 U3696 ( .A(n3005),  .B(n3287),  .C(n2452), .Y(w_mem_inst_n2051));
   AOI22X1 U3697 ( .A(block[84]),  .B(n3030),  .C(w_mem_inst_w_mem[52]),  .D(n3074), .Y(n3288));
   INVX1 U3698 ( .A(w_mem_inst_w_mem[84]), .Y(n3287));
   OAI21X1 U3699 ( .A(n3005),  .B(n3289),  .C(n2397), .Y(w_mem_inst_n2050));
   AOI22X1 U3700 ( .A(block[85]),  .B(n3030),  .C(w_mem_inst_w_mem[53]),  .D(n3074), .Y(n3290));
   INVX1 U3701 ( .A(w_mem_inst_w_mem[85]), .Y(n3289));
   OAI21X1 U3702 ( .A(n3005),  .B(n3291),  .C(n2794), .Y(w_mem_inst_n2049));
   AOI22X1 U3703 ( .A(block[86]),  .B(n3031),  .C(w_mem_inst_w_mem[54]),  .D(n3074), .Y(n3292));
   INVX1 U3704 ( .A(w_mem_inst_w_mem[86]), .Y(n3291));
   OAI21X1 U3705 ( .A(n3005),  .B(n3293),  .C(n2287), .Y(w_mem_inst_n2048));
   AOI22X1 U3706 ( .A(block[87]),  .B(n3031),  .C(w_mem_inst_w_mem[55]),  .D(n3074), .Y(n3294));
   INVX1 U3707 ( .A(w_mem_inst_w_mem[87]), .Y(n3293));
   OAI21X1 U3708 ( .A(n3005),  .B(n3295),  .C(n2335), .Y(w_mem_inst_n2047));
   AOI22X1 U3709 ( .A(block[88]),  .B(n3031),  .C(w_mem_inst_w_mem[56]),  .D(n3074), .Y(n3296));
   INVX1 U3710 ( .A(w_mem_inst_w_mem[88]), .Y(n3295));
   OAI21X1 U3711 ( .A(n3005),  .B(n3297),  .C(n2212), .Y(w_mem_inst_n2046));
   AOI22X1 U3712 ( .A(block[89]),  .B(n3031),  .C(w_mem_inst_w_mem[57]),  .D(n3074), .Y(n3298));
   INVX1 U3713 ( .A(w_mem_inst_w_mem[89]), .Y(n3297));
   OAI21X1 U3714 ( .A(n3005),  .B(n3299),  .C(n2238), .Y(w_mem_inst_n2045));
   AOI22X1 U3715 ( .A(block[90]),  .B(n3031),  .C(w_mem_inst_w_mem[58]),  .D(n3074), .Y(n3300));
   INVX1 U3716 ( .A(w_mem_inst_w_mem[90]), .Y(n3299));
   OAI21X1 U3717 ( .A(n3005),  .B(n3301),  .C(n2167), .Y(w_mem_inst_n2044));
   AOI22X1 U3718 ( .A(block[91]),  .B(n3031),  .C(w_mem_inst_w_mem[59]),  .D(n3074), .Y(n3302));
   INVX1 U3719 ( .A(w_mem_inst_w_mem[91]), .Y(n3301));
   OAI21X1 U3720 ( .A(n3004),  .B(n3303),  .C(n2437), .Y(w_mem_inst_n2043));
   AOI22X1 U3721 ( .A(block[92]),  .B(n3031),  .C(w_mem_inst_w_mem[60]),  .D(n3073), .Y(n3304));
   INVX1 U3722 ( .A(w_mem_inst_w_mem[92]), .Y(n3303));
   OAI21X1 U3723 ( .A(n3004),  .B(n3305),  .C(n2381), .Y(w_mem_inst_n2042));
   AOI22X1 U3724 ( .A(block[93]),  .B(n3031),  .C(w_mem_inst_w_mem[61]),  .D(n3073), .Y(n3306));
   INVX1 U3725 ( .A(w_mem_inst_w_mem[93]), .Y(n3305));
   OAI21X1 U3726 ( .A(n3004),  .B(n3307),  .C(n2182), .Y(w_mem_inst_n2041));
   AOI22X1 U3727 ( .A(block[94]),  .B(n3031),  .C(w_mem_inst_w_mem[62]),  .D(n3073), .Y(n3308));
   INVX1 U3728 ( .A(w_mem_inst_w_mem[94]), .Y(n3307));
   OAI21X1 U3729 ( .A(n3004),  .B(n3309),  .C(n2147), .Y(w_mem_inst_n2040));
   AOI22X1 U3730 ( .A(block[95]),  .B(n3031),  .C(w_mem_inst_w_mem[63]),  .D(n3073), .Y(n3310));
   INVX1 U3731 ( .A(w_mem_inst_w_mem[95]), .Y(n3309));
   OAI21X1 U3732 ( .A(n3004),  .B(n3311),  .C(n2884), .Y(w_mem_inst_n2039));
   AOI22X1 U3733 ( .A(block[96]),  .B(n3031),  .C(w_mem_inst_w_mem[64]),  .D(n3073), .Y(n3312));
   OAI21X1 U3734 ( .A(n3004),  .B(n3313),  .C(n2926), .Y(w_mem_inst_n2038));
   AOI22X1 U3735 ( .A(block[97]),  .B(n3031),  .C(w_mem_inst_w_mem[65]),  .D(n3073), .Y(n3314));
   OAI21X1 U3736 ( .A(n3004),  .B(n3315),  .C(n2762), .Y(w_mem_inst_n2037));
   AOI22X1 U3737 ( .A(block[98]),  .B(n3031),  .C(w_mem_inst_w_mem[66]),  .D(n3073), .Y(n3316));
   OAI21X1 U3738 ( .A(n3004),  .B(n3317),  .C(n2818), .Y(w_mem_inst_n2036));
   AOI22X1 U3739 ( .A(block[99]),  .B(n3032),  .C(w_mem_inst_w_mem[67]),  .D(n3073), .Y(n3318));
   OAI21X1 U3740 ( .A(n3004),  .B(n3319),  .C(n2698), .Y(w_mem_inst_n2035));
   AOI22X1 U3741 ( .A(block[100]),  .B(n3032),  .C(w_mem_inst_w_mem[68]),  .D(n3073), .Y(n3320));
   OAI21X1 U3742 ( .A(n3004),  .B(n3321),  .C(n2629), .Y(w_mem_inst_n2034));
   AOI22X1 U3743 ( .A(block[101]),  .B(n3032),  .C(w_mem_inst_w_mem[69]),  .D(n3073), .Y(n3322));
   OAI21X1 U3744 ( .A(n3004),  .B(n3323),  .C(n2579), .Y(w_mem_inst_n2033));
   AOI22X1 U3745 ( .A(block[102]),  .B(n3032),  .C(w_mem_inst_w_mem[70]),  .D(n3073), .Y(n3324));
   OAI21X1 U3746 ( .A(n3004),  .B(n3325),  .C(n2515), .Y(w_mem_inst_n2032));
   AOI22X1 U3747 ( .A(block[103]),  .B(n3032),  .C(w_mem_inst_w_mem[71]),  .D(n3073), .Y(n3326));
   OAI21X1 U3748 ( .A(n3003),  .B(n3327),  .C(n2918), .Y(w_mem_inst_n2031));
   AOI22X1 U3749 ( .A(block[104]),  .B(n3032),  .C(w_mem_inst_w_mem[72]),  .D(n3072), .Y(n3328));
   OAI21X1 U3750 ( .A(n3003),  .B(n3329),  .C(n2869), .Y(w_mem_inst_n2030));
   AOI22X1 U3751 ( .A(block[105]),  .B(n3032),  .C(w_mem_inst_w_mem[73]),  .D(n3072), .Y(n3330));
   OAI21X1 U3752 ( .A(n3003),  .B(n3331),  .C(n2746), .Y(w_mem_inst_n2029));
   AOI22X1 U3753 ( .A(block[106]),  .B(n3032),  .C(w_mem_inst_w_mem[74]),  .D(n3072), .Y(n3332));
   OAI21X1 U3754 ( .A(n3003),  .B(n3333),  .C(n2459), .Y(w_mem_inst_n2028));
   AOI22X1 U3755 ( .A(block[107]),  .B(n3032),  .C(w_mem_inst_w_mem[75]),  .D(n3072), .Y(n3334));
   OAI21X1 U3756 ( .A(n3003),  .B(n3335),  .C(n2404), .Y(w_mem_inst_n2027));
   AOI22X1 U3757 ( .A(block[108]),  .B(n3032),  .C(w_mem_inst_w_mem[76]),  .D(n3072), .Y(n3336));
   OAI21X1 U3758 ( .A(n3003),  .B(n3337),  .C(n2298), .Y(w_mem_inst_n2026));
   AOI22X1 U3759 ( .A(block[109]),  .B(n3032),  .C(w_mem_inst_w_mem[77]),  .D(n3072), .Y(n3338));
   OAI21X1 U3760 ( .A(n3003),  .B(n3339),  .C(n2348), .Y(w_mem_inst_n2025));
   AOI22X1 U3761 ( .A(block[110]),  .B(n3032),  .C(w_mem_inst_w_mem[78]),  .D(n3072), .Y(n3340));
   OAI21X1 U3762 ( .A(n3003),  .B(n3341),  .C(n2254), .Y(w_mem_inst_n2024));
   AOI22X1 U3763 ( .A(block[111]),  .B(n3032),  .C(w_mem_inst_w_mem[79]),  .D(n3072), .Y(n3342));
   OAI21X1 U3764 ( .A(n3003),  .B(n3343),  .C(n2798), .Y(w_mem_inst_n2023));
   AOI22X1 U3765 ( .A(block[112]),  .B(n3033),  .C(w_mem_inst_w_mem[80]),  .D(n3072), .Y(n3344));
   OAI21X1 U3766 ( .A(n3003),  .B(n3345),  .C(n2675), .Y(w_mem_inst_n2022));
   AOI22X1 U3767 ( .A(block[113]),  .B(n3033),  .C(w_mem_inst_w_mem[81]),  .D(n3072), .Y(n3346));
   OAI21X1 U3768 ( .A(n3003),  .B(n3347),  .C(n2613), .Y(w_mem_inst_n2021));
   AOI22X1 U3769 ( .A(block[114]),  .B(n3033),  .C(w_mem_inst_w_mem[82]),  .D(n3072), .Y(n3348));
   OAI21X1 U3770 ( .A(n3003),  .B(n3349),  .C(n2556), .Y(w_mem_inst_n2020));
   AOI22X1 U3771 ( .A(block[115]),  .B(n3033),  .C(w_mem_inst_w_mem[83]),  .D(n3072), .Y(n3350));
   OAI21X1 U3772 ( .A(n3002),  .B(n3351),  .C(n2902), .Y(w_mem_inst_n2019));
   AOI22X1 U3773 ( .A(block[116]),  .B(n3033),  .C(w_mem_inst_w_mem[84]),  .D(n3071), .Y(n3352));
   OAI21X1 U3774 ( .A(n3002),  .B(n3353),  .C(n2853), .Y(w_mem_inst_n2018));
   AOI22X1 U3775 ( .A(block[117]),  .B(n3033),  .C(w_mem_inst_w_mem[85]),  .D(n3071), .Y(n3354));
   OAI21X1 U3776 ( .A(n3002),  .B(n3355),  .C(n2731), .Y(w_mem_inst_n2017));
   AOI22X1 U3777 ( .A(block[118]),  .B(n3033),  .C(w_mem_inst_w_mem[86]),  .D(n3071), .Y(n3356));
   OAI21X1 U3778 ( .A(n3002),  .B(n3357),  .C(n2496), .Y(w_mem_inst_n2016));
   AOI22X1 U3779 ( .A(block[119]),  .B(n3033),  .C(w_mem_inst_w_mem[87]),  .D(n3071), .Y(n3358));
   OAI21X1 U3780 ( .A(n3002),  .B(n3359),  .C(n2443), .Y(w_mem_inst_n2015));
   AOI22X1 U3781 ( .A(block[120]),  .B(n3033),  .C(w_mem_inst_w_mem[88]),  .D(n3071), .Y(n3360));
   OAI21X1 U3782 ( .A(n3002),  .B(n3361),  .C(n2387), .Y(w_mem_inst_n2014));
   AOI22X1 U3783 ( .A(block[121]),  .B(n3033),  .C(w_mem_inst_w_mem[89]),  .D(n3071), .Y(n3362));
   OAI21X1 U3784 ( .A(n3002),  .B(n3363),  .C(n2332), .Y(w_mem_inst_n2013));
   AOI22X1 U3785 ( .A(block[122]),  .B(n3033),  .C(w_mem_inst_w_mem[90]),  .D(n3071), .Y(n3364));
   OAI21X1 U3786 ( .A(n3002),  .B(n3365),  .C(n2280), .Y(w_mem_inst_n2012));
   AOI22X1 U3787 ( .A(block[123]),  .B(n3033),  .C(w_mem_inst_w_mem[91]),  .D(n3071), .Y(n3366));
   OAI21X1 U3788 ( .A(n3002),  .B(n3367),  .C(n2236), .Y(w_mem_inst_n2011));
   AOI22X1 U3789 ( .A(block[124]),  .B(n3033),  .C(w_mem_inst_w_mem[92]),  .D(n3071), .Y(n3368));
   OAI21X1 U3790 ( .A(n3002),  .B(n3369),  .C(n2204), .Y(w_mem_inst_n2010));
   AOI22X1 U3791 ( .A(block[125]),  .B(n3034),  .C(w_mem_inst_w_mem[93]),  .D(n3071), .Y(n3370));
   OAI21X1 U3792 ( .A(n3002),  .B(n3371),  .C(n2161), .Y(w_mem_inst_n2009));
   AOI22X1 U3793 ( .A(block[126]),  .B(n3034),  .C(w_mem_inst_w_mem[94]),  .D(n3071), .Y(n3372));
   OAI21X1 U3794 ( .A(n3002),  .B(n3373),  .C(n2178), .Y(w_mem_inst_n2008));
   AOI22X1 U3795 ( .A(block[127]),  .B(n3034),  .C(w_mem_inst_w_mem[95]),  .D(n3071), .Y(n3374));
   OAI21X1 U3796 ( .A(n3001),  .B(n3375),  .C(n2933), .Y(w_mem_inst_n2007));
   AOI22X1 U3797 ( .A(block[128]),  .B(n3034),  .C(w_mem_inst_w_mem[96]),  .D(n3070), .Y(n3376));
   INVX1 U3798 ( .A(w_mem_inst_w_mem[128]), .Y(n3375));
   OAI21X1 U3799 ( .A(n3001),  .B(n3377),  .C(n2875), .Y(w_mem_inst_n2006));
   AOI22X1 U3800 ( .A(block[129]),  .B(n3034),  .C(w_mem_inst_w_mem[97]),  .D(n3070), .Y(n3378));
   INVX1 U3801 ( .A(w_mem_inst_w_mem[129]), .Y(n3377));
   OAI21X1 U3802 ( .A(n3001),  .B(n3379),  .C(n2825), .Y(w_mem_inst_n2005));
   AOI22X1 U3803 ( .A(block[130]),  .B(n3034),  .C(w_mem_inst_w_mem[98]),  .D(n3070), .Y(n3380));
   OAI21X1 U3804 ( .A(n3001),  .B(n3381),  .C(n2753), .Y(w_mem_inst_n2004));
   AOI22X1 U3805 ( .A(block[131]),  .B(n3034),  .C(w_mem_inst_w_mem[99]),  .D(n3070), .Y(n3382));
   OAI21X1 U3806 ( .A(n3001),  .B(n3383),  .C(n2635), .Y(w_mem_inst_n2003));
   AOI22X1 U3807 ( .A(block[132]),  .B(n3034),  .C(w_mem_inst_w_mem[100]),  .D(n3070), .Y(n3384));
   OAI21X1 U3808 ( .A(n3001),  .B(n3385),  .C(n2691), .Y(w_mem_inst_n2002));
   AOI22X1 U3809 ( .A(block[133]),  .B(n3034),  .C(w_mem_inst_w_mem[101]),  .D(n3070), .Y(n3386));
   OAI21X1 U3810 ( .A(n3001),  .B(n3387),  .C(n2521), .Y(w_mem_inst_n2001));
   AOI22X1 U3811 ( .A(block[134]),  .B(n3034),  .C(w_mem_inst_w_mem[102]),  .D(n3070), .Y(n3388));
   OAI21X1 U3812 ( .A(n3001),  .B(n3389),  .C(n2572), .Y(w_mem_inst_n2000));
   AOI22X1 U3813 ( .A(block[135]),  .B(n3034),  .C(w_mem_inst_w_mem[103]),  .D(n3070), .Y(n3390));
   OAI21X1 U3814 ( .A(n3001),  .B(n3391),  .C(n2467), .Y(w_mem_inst_n1999));
   AOI22X1 U3815 ( .A(block[136]),  .B(n3034),  .C(w_mem_inst_w_mem[104]),  .D(n3070), .Y(n3392));
   OAI21X1 U3816 ( .A(n3001),  .B(n3393),  .C(n2409), .Y(w_mem_inst_n1998));
   AOI22X1 U3817 ( .A(block[137]),  .B(n3034),  .C(w_mem_inst_w_mem[105]),  .D(n3070), .Y(n3394));
   OAI21X1 U3818 ( .A(n3001),  .B(n3395),  .C(n2355), .Y(w_mem_inst_n1997));
   AOI22X1 U3819 ( .A(block[138]),  .B(n3035),  .C(w_mem_inst_w_mem[106]),  .D(n3070), .Y(n3396));
   INVX1 U3820 ( .A(w_mem_inst_w_mem[138]), .Y(n3395));
   OAI21X1 U3821 ( .A(n3001),  .B(n3397),  .C(n2302), .Y(w_mem_inst_n1996));
   AOI22X1 U3822 ( .A(block[139]),  .B(n3035),  .C(w_mem_inst_w_mem[107]),  .D(n3070), .Y(n3398));
   INVX1 U3823 ( .A(w_mem_inst_w_mem[139]), .Y(n3397));
   OAI21X1 U3824 ( .A(n3000),  .B(n3399),  .C(n2907), .Y(w_mem_inst_n1995));
   AOI22X1 U3825 ( .A(block[140]),  .B(n3035),  .C(w_mem_inst_w_mem[108]),  .D(n3069), .Y(n3400));
   INVX1 U3826 ( .A(w_mem_inst_w_mem[140]), .Y(n3399));
   OAI21X1 U3827 ( .A(n3000),  .B(n3401),  .C(n2857), .Y(w_mem_inst_n1994));
   AOI22X1 U3828 ( .A(block[141]),  .B(n3035),  .C(w_mem_inst_w_mem[109]),  .D(n3069), .Y(n3402));
   INVX1 U3829 ( .A(w_mem_inst_w_mem[141]), .Y(n3401));
   OAI21X1 U3830 ( .A(n3000),  .B(n3403),  .C(n2802), .Y(w_mem_inst_n1993));
   AOI22X1 U3831 ( .A(block[142]),  .B(n3035),  .C(w_mem_inst_w_mem[110]),  .D(n3069), .Y(n3404));
   INVX1 U3832 ( .A(w_mem_inst_w_mem[142]), .Y(n3403));
   OAI21X1 U3833 ( .A(n3000),  .B(n3405),  .C(n2737), .Y(w_mem_inst_n1992));
   AOI22X1 U3834 ( .A(block[143]),  .B(n3035),  .C(w_mem_inst_w_mem[111]),  .D(n3069), .Y(n3406));
   INVX1 U3835 ( .A(w_mem_inst_w_mem[143]), .Y(n3405));
   OAI21X1 U3836 ( .A(n3000),  .B(n3407),  .C(n2680), .Y(w_mem_inst_n1991));
   AOI22X1 U3837 ( .A(block[144]),  .B(n3035),  .C(w_mem_inst_w_mem[112]),  .D(n3069), .Y(n3408));
   INVX1 U3838 ( .A(w_mem_inst_w_mem[144]), .Y(n3407));
   OAI21X1 U3839 ( .A(n3000),  .B(n3409),  .C(n2618), .Y(w_mem_inst_n1990));
   AOI22X1 U3840 ( .A(block[145]),  .B(n3035),  .C(w_mem_inst_w_mem[113]),  .D(n3069), .Y(n3410));
   INVX1 U3841 ( .A(w_mem_inst_w_mem[145]), .Y(n3409));
   OAI21X1 U3842 ( .A(n3000),  .B(n3411),  .C(n2561), .Y(w_mem_inst_n1989));
   AOI22X1 U3843 ( .A(block[146]),  .B(n3035),  .C(w_mem_inst_w_mem[114]),  .D(n3069), .Y(n3412));
   INVX1 U3844 ( .A(w_mem_inst_w_mem[146]), .Y(n3411));
   OAI21X1 U3845 ( .A(n3000),  .B(n3413),  .C(n2504), .Y(w_mem_inst_n1988));
   AOI22X1 U3846 ( .A(block[147]),  .B(n3035),  .C(w_mem_inst_w_mem[115]),  .D(n3069), .Y(n3414));
   INVX1 U3847 ( .A(w_mem_inst_w_mem[147]), .Y(n3413));
   OAI21X1 U3848 ( .A(n3000),  .B(n3415),  .C(n2451), .Y(w_mem_inst_n1987));
   AOI22X1 U3849 ( .A(block[148]),  .B(n3035),  .C(w_mem_inst_w_mem[116]),  .D(n3069), .Y(n3416));
   INVX1 U3850 ( .A(w_mem_inst_w_mem[148]), .Y(n3415));
   OAI21X1 U3851 ( .A(n3000),  .B(n3417),  .C(n2396), .Y(w_mem_inst_n1986));
   AOI22X1 U3852 ( .A(block[149]),  .B(n3035),  .C(w_mem_inst_w_mem[117]),  .D(n3069), .Y(n3418));
   INVX1 U3853 ( .A(w_mem_inst_w_mem[149]), .Y(n3417));
   OAI21X1 U3854 ( .A(n3000),  .B(n3419),  .C(n2246), .Y(w_mem_inst_n1985));
   AOI22X1 U3855 ( .A(block[150]),  .B(n3035),  .C(w_mem_inst_w_mem[118]),  .D(n3069), .Y(n3420));
   INVX1 U3856 ( .A(w_mem_inst_w_mem[150]), .Y(n3419));
   OAI21X1 U3857 ( .A(n3000),  .B(n3421),  .C(n2339), .Y(w_mem_inst_n1984));
   AOI22X1 U3858 ( .A(block[151]),  .B(n3036),  .C(w_mem_inst_w_mem[119]),  .D(n3069), .Y(n3422));
   OAI21X1 U3859 ( .A(n2999),  .B(n3423),  .C(n2667), .Y(w_mem_inst_n1983));
   AOI22X1 U3860 ( .A(block[152]),  .B(n3036),  .C(w_mem_inst_w_mem[120]),  .D(n3068), .Y(n3424));
   OAI21X1 U3861 ( .A(n2999),  .B(n3425),  .C(n2603), .Y(w_mem_inst_n1982));
   AOI22X1 U3862 ( .A(block[153]),  .B(n3036),  .C(w_mem_inst_w_mem[121]),  .D(n3068), .Y(n3426));
   OAI21X1 U3863 ( .A(n2999),  .B(n3427),  .C(n2547), .Y(w_mem_inst_n1981));
   AOI22X1 U3864 ( .A(block[154]),  .B(n3036),  .C(w_mem_inst_w_mem[122]),  .D(n3068), .Y(n3428));
   OAI21X1 U3865 ( .A(n2999),  .B(n3429),  .C(n2489), .Y(w_mem_inst_n1980));
   AOI22X1 U3866 ( .A(block[155]),  .B(n3036),  .C(w_mem_inst_w_mem[123]),  .D(n3068), .Y(n3430));
   OAI21X1 U3867 ( .A(n2999),  .B(n3431),  .C(n2436), .Y(w_mem_inst_n1979));
   AOI22X1 U3868 ( .A(block[156]),  .B(n3036),  .C(w_mem_inst_w_mem[124]),  .D(n3068), .Y(n3432));
   OAI21X1 U3869 ( .A(n2999),  .B(n3433),  .C(n2380), .Y(w_mem_inst_n1978));
   AOI22X1 U3870 ( .A(block[157]),  .B(n3036),  .C(w_mem_inst_w_mem[125]),  .D(n3068), .Y(n3434));
   OAI21X1 U3871 ( .A(n2999),  .B(n3435),  .C(n2273), .Y(w_mem_inst_n1977));
   AOI22X1 U3872 ( .A(block[158]),  .B(n3036),  .C(w_mem_inst_w_mem[126]),  .D(n3068), .Y(n3436));
   OAI21X1 U3873 ( .A(n2999),  .B(n3437),  .C(n2230), .Y(w_mem_inst_n1976));
   AOI22X1 U3874 ( .A(block[159]),  .B(n3036),  .C(w_mem_inst_w_mem[127]),  .D(n3068), .Y(n3438));
   OAI21X1 U3875 ( .A(n2999),  .B(n3439),  .C(n2883), .Y(w_mem_inst_n1975));
   AOI22X1 U3876 ( .A(block[160]),  .B(n3036),  .C(w_mem_inst_w_mem[128]),  .D(n3068), .Y(n3440));
   OAI21X1 U3877 ( .A(n2999),  .B(n3441),  .C(n2925), .Y(w_mem_inst_n1974));
   AOI22X1 U3878 ( .A(block[161]),  .B(n3036),  .C(w_mem_inst_w_mem[129]),  .D(n3068), .Y(n3442));
   OAI21X1 U3879 ( .A(n2999),  .B(n3443),  .C(n2761), .Y(w_mem_inst_n1973));
   AOI22X1 U3880 ( .A(block[162]),  .B(n3036),  .C(w_mem_inst_w_mem[130]),  .D(n3068), .Y(n3444));
   OAI21X1 U3881 ( .A(n2999),  .B(n3445),  .C(n2817), .Y(w_mem_inst_n1972));
   AOI22X1 U3882 ( .A(block[163]),  .B(n3018),  .C(w_mem_inst_w_mem[131]),  .D(n3068), .Y(n3446));
   OAI21X1 U3883 ( .A(n2998),  .B(n3447),  .C(n2919), .Y(w_mem_inst_n1971));
   AOI22X1 U3884 ( .A(block[164]),  .B(n3013),  .C(w_mem_inst_w_mem[132]),  .D(n3067), .Y(n3448));
   OAI21X1 U3885 ( .A(n2998),  .B(n3449),  .C(n2811), .Y(w_mem_inst_n1970));
   AOI22X1 U3886 ( .A(block[165]),  .B(n3013),  .C(w_mem_inst_w_mem[133]),  .D(n3067), .Y(n3450));
   OAI21X1 U3887 ( .A(n2998),  .B(n3451),  .C(n2747), .Y(w_mem_inst_n1969));
   AOI22X1 U3888 ( .A(block[166]),  .B(n3013),  .C(w_mem_inst_w_mem[134]),  .D(n3067), .Y(n3452));
   OAI21X1 U3889 ( .A(n2998),  .B(n3453),  .C(n2686), .Y(w_mem_inst_n1968));
   AOI22X1 U3890 ( .A(block[167]),  .B(n3013),  .C(w_mem_inst_w_mem[135]),  .D(n3067), .Y(n3454));
   OAI21X1 U3891 ( .A(n2998),  .B(n3455),  .C(n2622), .Y(w_mem_inst_n1967));
   AOI22X1 U3892 ( .A(block[168]),  .B(n3013),  .C(w_mem_inst_w_mem[136]),  .D(n3067), .Y(n3456));
   OAI21X1 U3893 ( .A(n2998),  .B(n3457),  .C(n2567), .Y(w_mem_inst_n1966));
   AOI22X1 U3894 ( .A(block[169]),  .B(n3013),  .C(w_mem_inst_w_mem[137]),  .D(n3067), .Y(n3458));
   OAI21X1 U3895 ( .A(n2998),  .B(n3459),  .C(n2508), .Y(w_mem_inst_n1965));
   AOI22X1 U3896 ( .A(block[170]),  .B(n3013),  .C(w_mem_inst_w_mem[138]),  .D(n3067), .Y(n3460));
   OAI21X1 U3897 ( .A(n2998),  .B(n3461),  .C(n2458), .Y(w_mem_inst_n1964));
   AOI22X1 U3898 ( .A(block[171]),  .B(n3013),  .C(w_mem_inst_w_mem[139]),  .D(n3067), .Y(n3462));
   OAI21X1 U3899 ( .A(n2998),  .B(n3463),  .C(n2403), .Y(w_mem_inst_n1963));
   AOI22X1 U3900 ( .A(block[172]),  .B(n3013),  .C(w_mem_inst_w_mem[140]),  .D(n3067), .Y(n3464));
   OAI21X1 U3901 ( .A(n2998),  .B(n3465),  .C(n2350), .Y(w_mem_inst_n1962));
   AOI22X1 U3902 ( .A(block[173]),  .B(n3013),  .C(w_mem_inst_w_mem[141]),  .D(n3067), .Y(n3466));
   OAI21X1 U3903 ( .A(n2998),  .B(n3467),  .C(n2296), .Y(w_mem_inst_n1961));
   AOI22X1 U3904 ( .A(block[174]),  .B(n3013),  .C(w_mem_inst_w_mem[142]),  .D(n3067), .Y(n3468));
   OAI21X1 U3905 ( .A(n2998),  .B(n3469),  .C(n2253), .Y(w_mem_inst_n1960));
   AOI22X1 U3906 ( .A(block[175]),  .B(n3013),  .C(w_mem_inst_w_mem[143]),  .D(n3067), .Y(n3470));
   OAI21X1 U3907 ( .A(n2997),  .B(n3471),  .C(n2904), .Y(w_mem_inst_n1959));
   AOI22X1 U3908 ( .A(block[176]),  .B(n3014),  .C(w_mem_inst_w_mem[144]),  .D(n3066), .Y(n3472));
   OAI21X1 U3909 ( .A(n2997),  .B(n3473),  .C(n2854), .Y(w_mem_inst_n1958));
   AOI22X1 U3910 ( .A(block[177]),  .B(n3014),  .C(w_mem_inst_w_mem[145]),  .D(n3066), .Y(n3474));
   OAI21X1 U3911 ( .A(n2997),  .B(n3475),  .C(n2796), .Y(w_mem_inst_n1957));
   AOI22X1 U3912 ( .A(block[178]),  .B(n3014),  .C(w_mem_inst_w_mem[146]),  .D(n3066), .Y(n3476));
   OAI21X1 U3913 ( .A(n2997),  .B(n3477),  .C(n2732), .Y(w_mem_inst_n1956));
   AOI22X1 U3914 ( .A(block[179]),  .B(n3014),  .C(w_mem_inst_w_mem[147]),  .D(n3066), .Y(n3478));
   OAI21X1 U3915 ( .A(n2997),  .B(n3479),  .C(n2670), .Y(w_mem_inst_n1955));
   AOI22X1 U3916 ( .A(block[180]),  .B(n3014),  .C(w_mem_inst_w_mem[148]),  .D(n3066), .Y(n3480));
   OAI21X1 U3917 ( .A(n2997),  .B(n3481),  .C(n2606), .Y(w_mem_inst_n1954));
   AOI22X1 U3918 ( .A(block[181]),  .B(n3014),  .C(w_mem_inst_w_mem[149]),  .D(n3066), .Y(n3482));
   OAI21X1 U3919 ( .A(n2997),  .B(n3483),  .C(n2551), .Y(w_mem_inst_n1953));
   AOI22X1 U3920 ( .A(block[182]),  .B(n3014),  .C(w_mem_inst_w_mem[150]),  .D(n3066), .Y(n3484));
   OAI21X1 U3921 ( .A(n2997),  .B(n3485),  .C(n2495), .Y(w_mem_inst_n1952));
   AOI22X1 U3922 ( .A(block[183]),  .B(n3014),  .C(w_mem_inst_w_mem[151]),  .D(n3066), .Y(n3486));
   OAI21X1 U3923 ( .A(n2997),  .B(n3487),  .C(n2442), .Y(w_mem_inst_n1951));
   AOI22X1 U3924 ( .A(block[184]),  .B(n3014),  .C(w_mem_inst_w_mem[152]),  .D(n3066), .Y(n3488));
   OAI21X1 U3925 ( .A(n2997),  .B(n3489),  .C(n2386), .Y(w_mem_inst_n1950));
   AOI22X1 U3926 ( .A(block[185]),  .B(n3014),  .C(w_mem_inst_w_mem[153]),  .D(n3066), .Y(n3490));
   OAI21X1 U3927 ( .A(n2997),  .B(n3491),  .C(n2331), .Y(w_mem_inst_n1949));
   AOI22X1 U3928 ( .A(block[186]),  .B(n3014),  .C(w_mem_inst_w_mem[154]),  .D(n3066), .Y(n3492));
   OAI21X1 U3929 ( .A(n2997),  .B(n3493),  .C(n2279), .Y(w_mem_inst_n1948));
   AOI22X1 U3930 ( .A(block[187]),  .B(n3014),  .C(w_mem_inst_w_mem[155]),  .D(n3066), .Y(n3494));
   OAI21X1 U3931 ( .A(n2996),  .B(n3495),  .C(n2235), .Y(w_mem_inst_n1947));
   AOI22X1 U3932 ( .A(block[188]),  .B(n3014),  .C(w_mem_inst_w_mem[156]),  .D(n3065), .Y(n3496));
   OAI21X1 U3933 ( .A(n2996),  .B(n3497),  .C(n2325), .Y(w_mem_inst_n1946));
   AOI22X1 U3934 ( .A(block[189]),  .B(n3015),  .C(w_mem_inst_w_mem[157]),  .D(n3065), .Y(n3498));
   OAI21X1 U3935 ( .A(n2996),  .B(n3499),  .C(n2201), .Y(w_mem_inst_n1945));
   AOI22X1 U3936 ( .A(block[190]),  .B(n3015),  .C(w_mem_inst_w_mem[158]),  .D(n3065), .Y(n3500));
   OAI21X1 U3937 ( .A(n2996),  .B(n3501),  .C(n2271), .Y(w_mem_inst_n1944));
   AOI22X1 U3938 ( .A(block[191]),  .B(n3015),  .C(w_mem_inst_w_mem[159]),  .D(n3065), .Y(n3502));
   OAI21X1 U3939 ( .A(n2996),  .B(n3503),  .C(n2932), .Y(w_mem_inst_n1943));
   AOI22X1 U3940 ( .A(block[192]),  .B(n3015),  .C(w_mem_inst_w_mem[160]),  .D(n3065), .Y(n3504));
   OAI21X1 U3941 ( .A(n2996),  .B(n3505),  .C(n2874), .Y(w_mem_inst_n1942));
   AOI22X1 U3942 ( .A(block[193]),  .B(n3015),  .C(w_mem_inst_w_mem[161]),  .D(n3065), .Y(n3506));
   OAI21X1 U3943 ( .A(n2996),  .B(n3507),  .C(n2824), .Y(w_mem_inst_n1941));
   AOI22X1 U3944 ( .A(block[194]),  .B(n3015),  .C(w_mem_inst_w_mem[162]),  .D(n3065), .Y(n3508));
   OAI21X1 U3945 ( .A(n2996),  .B(n3509),  .C(n2752), .Y(w_mem_inst_n1940));
   AOI22X1 U3946 ( .A(block[195]),  .B(n3015),  .C(w_mem_inst_w_mem[163]),  .D(n3065), .Y(n3510));
   OAI21X1 U3947 ( .A(n2996),  .B(n3511),  .C(n2697), .Y(w_mem_inst_n1939));
   AOI22X1 U3948 ( .A(block[196]),  .B(n3015),  .C(w_mem_inst_w_mem[164]),  .D(n3065), .Y(n3512));
   OAI21X1 U3949 ( .A(n2996),  .B(n3513),  .C(n2628), .Y(w_mem_inst_n1938));
   AOI22X1 U3950 ( .A(block[197]),  .B(n3015),  .C(w_mem_inst_w_mem[165]),  .D(n3065), .Y(n3514));
   OAI21X1 U3951 ( .A(n2996),  .B(n3515),  .C(n2578), .Y(w_mem_inst_n1937));
   AOI22X1 U3952 ( .A(block[198]),  .B(n3015),  .C(w_mem_inst_w_mem[166]),  .D(n3065), .Y(n3516));
   OAI21X1 U3953 ( .A(n2996),  .B(n3517),  .C(n2514), .Y(w_mem_inst_n1936));
   AOI22X1 U3954 ( .A(block[199]),  .B(n3015),  .C(w_mem_inst_w_mem[167]),  .D(n3065), .Y(n3518));
   OAI21X1 U3955 ( .A(n2995),  .B(n3519),  .C(n2466), .Y(w_mem_inst_n1935));
   AOI22X1 U3956 ( .A(block[200]),  .B(n3015),  .C(w_mem_inst_w_mem[168]),  .D(n3064), .Y(n3520));
   OAI21X1 U3957 ( .A(n2995),  .B(n3521),  .C(n2408), .Y(w_mem_inst_n1934));
   AOI22X1 U3958 ( .A(block[201]),  .B(n3015),  .C(w_mem_inst_w_mem[169]),  .D(n3064), .Y(n3522));
   OAI21X1 U3959 ( .A(n2995),  .B(n3523),  .C(n2912), .Y(w_mem_inst_n1933));
   AOI22X1 U3960 ( .A(block[202]),  .B(n3016),  .C(w_mem_inst_w_mem[170]),  .D(n3064), .Y(n3524));
   OAI21X1 U3961 ( .A(n2995),  .B(n3525),  .C(n2863), .Y(w_mem_inst_n1932));
   AOI22X1 U3962 ( .A(block[203]),  .B(n3016),  .C(w_mem_inst_w_mem[171]),  .D(n3064), .Y(n3526));
   OAI21X1 U3963 ( .A(n2995),  .B(n3527),  .C(n2806), .Y(w_mem_inst_n1931));
   AOI22X1 U3964 ( .A(block[204]),  .B(n3016),  .C(w_mem_inst_w_mem[172]),  .D(n3064), .Y(n3528));
   OAI21X1 U3965 ( .A(n2995),  .B(n3529),  .C(n2741), .Y(w_mem_inst_n1930));
   AOI22X1 U3966 ( .A(block[205]),  .B(n3016),  .C(w_mem_inst_w_mem[173]),  .D(n3064), .Y(n3530));
   OAI21X1 U3967 ( .A(n2995),  .B(n3531),  .C(n2682), .Y(w_mem_inst_n1929));
   AOI22X1 U3968 ( .A(block[206]),  .B(n3016),  .C(w_mem_inst_w_mem[174]),  .D(n3064), .Y(n3532));
   OAI21X1 U3969 ( .A(n2995),  .B(n3533),  .C(n2620), .Y(w_mem_inst_n1928));
   AOI22X1 U3970 ( .A(block[207]),  .B(n3016),  .C(w_mem_inst_w_mem[175]),  .D(n3064), .Y(n3534));
   OAI21X1 U3971 ( .A(n2995),  .B(n3535),  .C(n2564), .Y(w_mem_inst_n1927));
   AOI22X1 U3972 ( .A(block[208]),  .B(n3016),  .C(w_mem_inst_w_mem[176]),  .D(n3064), .Y(n3536));
   OAI21X1 U3973 ( .A(n2995),  .B(n3537),  .C(n2506), .Y(w_mem_inst_n1926));
   AOI22X1 U3974 ( .A(block[209]),  .B(n3016),  .C(w_mem_inst_w_mem[177]),  .D(n3064), .Y(n3538));
   OAI21X1 U3975 ( .A(n2995),  .B(n3539),  .C(n2343), .Y(w_mem_inst_n1925));
   AOI22X1 U3976 ( .A(block[210]),  .B(n3016),  .C(w_mem_inst_w_mem[178]),  .D(n3064), .Y(n3540));
   OAI21X1 U3977 ( .A(n2995),  .B(n3541),  .C(n2289), .Y(w_mem_inst_n1924));
   AOI22X1 U3978 ( .A(block[211]),  .B(n3016),  .C(w_mem_inst_w_mem[179]),  .D(n3064), .Y(n3542));
   OAI21X1 U3979 ( .A(n2994),  .B(n3543),  .C(n2450), .Y(w_mem_inst_n1923));
   AOI22X1 U3980 ( .A(block[212]),  .B(n3016),  .C(w_mem_inst_w_mem[180]),  .D(n3063), .Y(n3544));
   OAI21X1 U3981 ( .A(n2994),  .B(n3545),  .C(n2395), .Y(w_mem_inst_n1922));
   AOI22X1 U3982 ( .A(block[213]),  .B(n3016),  .C(w_mem_inst_w_mem[181]),  .D(n3063), .Y(n3546));
   OAI21X1 U3983 ( .A(n2994),  .B(n3547),  .C(n2245), .Y(w_mem_inst_n1921));
   AOI22X1 U3984 ( .A(block[214]),  .B(n3016),  .C(w_mem_inst_w_mem[182]),  .D(n3063), .Y(n3548));
   OAI21X1 U3985 ( .A(n2994),  .B(n3549),  .C(n2668), .Y(w_mem_inst_n1920));
   AOI22X1 U3986 ( .A(block[215]),  .B(n3029),  .C(w_mem_inst_w_mem[183]),  .D(n3063), .Y(n3550));
   OAI21X1 U3987 ( .A(n2994),  .B(n3551),  .C(n2604), .Y(w_mem_inst_n1919));
   AOI22X1 U3988 ( .A(block[216]),  .B(n3027),  .C(w_mem_inst_w_mem[184]),  .D(n3063), .Y(n3552));
   OAI21X1 U3989 ( .A(n2994),  .B(n3553),  .C(n2549), .Y(w_mem_inst_n1918));
   AOI22X1 U3990 ( .A(block[217]),  .B(n3038),  .C(w_mem_inst_w_mem[185]),  .D(n3063), .Y(n3554));
   OAI21X1 U3991 ( .A(n2994),  .B(n3555),  .C(n2490), .Y(w_mem_inst_n1917));
   AOI22X1 U3992 ( .A(block[218]),  .B(n3034),  .C(w_mem_inst_w_mem[186]),  .D(n3063), .Y(n3556));
   OAI21X1 U3993 ( .A(n2994),  .B(n3557),  .C(n2329), .Y(w_mem_inst_n1916));
   AOI22X1 U3994 ( .A(block[219]),  .B(n3018),  .C(w_mem_inst_w_mem[187]),  .D(n3063), .Y(n3558));
   OAI21X1 U3995 ( .A(n2994),  .B(n3559),  .C(n2277), .Y(w_mem_inst_n1915));
   AOI22X1 U3996 ( .A(block[220]),  .B(n3037),  .C(w_mem_inst_w_mem[188]),  .D(n3063), .Y(n3560));
   OAI21X1 U3997 ( .A(n2994),  .B(n3561),  .C(n2203), .Y(w_mem_inst_n1914));
   AOI22X1 U3998 ( .A(block[221]),  .B(n3039),  .C(w_mem_inst_w_mem[189]),  .D(n3063), .Y(n3562));
   OAI21X1 U3999 ( .A(n2994),  .B(n3563),  .C(n2181), .Y(w_mem_inst_n1913));
   AOI22X1 U4000 ( .A(block[222]),  .B(n3048),  .C(w_mem_inst_w_mem[190]),  .D(n3063), .Y(n3564));
   OAI21X1 U4001 ( .A(n2994),  .B(n3565),  .C(n2159), .Y(w_mem_inst_n1912));
   AOI22X1 U4002 ( .A(block[223]),  .B(n3041),  .C(w_mem_inst_w_mem[191]),  .D(n3063), .Y(n3566));
   OAI21X1 U4003 ( .A(n2993),  .B(n3567),  .C(n2882), .Y(w_mem_inst_n1911));
   AOI22X1 U4004 ( .A(block[224]),  .B(n3050),  .C(w_mem_inst_w_mem[192]),  .D(n3062), .Y(n3568));
   OAI21X1 U4005 ( .A(n2993),  .B(n3569),  .C(n2924), .Y(w_mem_inst_n1910));
   AOI22X1 U4006 ( .A(block[225]),  .B(n3043),  .C(w_mem_inst_w_mem[193]),  .D(n3062), .Y(n3570));
   OAI21X1 U4007 ( .A(n2993),  .B(n3571),  .C(n2760), .Y(w_mem_inst_n1909));
   AOI22X1 U4008 ( .A(block[226]),  .B(n3045),  .C(w_mem_inst_w_mem[194]),  .D(n3062), .Y(n3572));
   OAI21X1 U4009 ( .A(n2993),  .B(n3573),  .C(n2816), .Y(w_mem_inst_n1908));
   AOI22X1 U4010 ( .A(block[227]),  .B(n3047),  .C(w_mem_inst_w_mem[195]),  .D(n3062), .Y(n3574));
   OAI21X1 U4011 ( .A(n2993),  .B(n3575),  .C(n2634), .Y(w_mem_inst_n1907));
   AOI22X1 U4012 ( .A(block[228]),  .B(n3017),  .C(w_mem_inst_w_mem[196]),  .D(n3062), .Y(n3576));
   OAI21X1 U4013 ( .A(n2993),  .B(n3577),  .C(n2690), .Y(w_mem_inst_n1906));
   AOI22X1 U4014 ( .A(block[229]),  .B(n3017),  .C(w_mem_inst_w_mem[197]),  .D(n3062), .Y(n3578));
   OAI21X1 U4015 ( .A(n2993),  .B(n3579),  .C(n2520), .Y(w_mem_inst_n1905));
   AOI22X1 U4016 ( .A(block[230]),  .B(n3017),  .C(w_mem_inst_w_mem[198]),  .D(n3062), .Y(n3580));
   OAI21X1 U4017 ( .A(n2993),  .B(n3581),  .C(n2571), .Y(w_mem_inst_n1904));
   AOI22X1 U4018 ( .A(block[231]),  .B(n3017),  .C(w_mem_inst_w_mem[199]),  .D(n3062), .Y(n3582));
   OAI21X1 U4019 ( .A(n2993),  .B(n3583),  .C(n2412), .Y(w_mem_inst_n1903));
   AOI22X1 U4020 ( .A(block[232]),  .B(n3017),  .C(w_mem_inst_w_mem[200]),  .D(n3062), .Y(n3584));
   OAI21X1 U4021 ( .A(n2993),  .B(n3585),  .C(n2461), .Y(w_mem_inst_n1902));
   AOI22X1 U4022 ( .A(block[233]),  .B(n3017),  .C(w_mem_inst_w_mem[201]),  .D(n3062), .Y(n3586));
   OAI21X1 U4023 ( .A(n2993),  .B(n3587),  .C(n2354), .Y(w_mem_inst_n1901));
   AOI22X1 U4024 ( .A(block[234]),  .B(n3017),  .C(w_mem_inst_w_mem[202]),  .D(n3062), .Y(n3588));
   OAI21X1 U4025 ( .A(n2993),  .B(n3589),  .C(n2301), .Y(w_mem_inst_n1900));
   AOI22X1 U4026 ( .A(block[235]),  .B(n3017),  .C(w_mem_inst_w_mem[203]),  .D(n3062), .Y(n3590));
   OAI21X1 U4027 ( .A(n2992),  .B(n3591),  .C(n2906), .Y(w_mem_inst_n1899));
   AOI22X1 U4028 ( .A(block[236]),  .B(n3017),  .C(w_mem_inst_w_mem[204]),  .D(n3061), .Y(n3592));
   OAI21X1 U4029 ( .A(n2992),  .B(n3593),  .C(n2856), .Y(w_mem_inst_n1898));
   AOI22X1 U4030 ( .A(block[237]),  .B(n3017),  .C(w_mem_inst_w_mem[205]),  .D(n3061), .Y(n3594));
   OAI21X1 U4031 ( .A(n2992),  .B(n3595),  .C(n2801), .Y(w_mem_inst_n1897));
   AOI22X1 U4032 ( .A(block[238]),  .B(n3017),  .C(w_mem_inst_w_mem[206]),  .D(n3061), .Y(n3596));
   OAI21X1 U4033 ( .A(n2992),  .B(n3597),  .C(n2736), .Y(w_mem_inst_n1896));
   AOI22X1 U4034 ( .A(block[239]),  .B(n3017),  .C(w_mem_inst_w_mem[207]),  .D(n3061), .Y(n3598));
   OAI21X1 U4035 ( .A(n2992),  .B(n3599),  .C(n2251), .Y(w_mem_inst_n1895));
   AOI22X1 U4036 ( .A(block[240]),  .B(n3017),  .C(w_mem_inst_w_mem[208]),  .D(n3061), .Y(n3600));
   OAI21X1 U4037 ( .A(n2992),  .B(n3601),  .C(n2674), .Y(w_mem_inst_n1894));
   AOI22X1 U4038 ( .A(block[241]),  .B(n3018),  .C(w_mem_inst_w_mem[209]),  .D(n3061), .Y(n3602));
   OAI21X1 U4039 ( .A(n2992),  .B(n3603),  .C(n2612), .Y(w_mem_inst_n1893));
   AOI22X1 U4040 ( .A(block[242]),  .B(n3018),  .C(w_mem_inst_w_mem[210]),  .D(n3061), .Y(n3604));
   OAI21X1 U4041 ( .A(n2992),  .B(n3605),  .C(n2555), .Y(w_mem_inst_n1892));
   AOI22X1 U4042 ( .A(block[243]),  .B(n3018),  .C(w_mem_inst_w_mem[211]),  .D(n3061), .Y(n3606));
   OAI21X1 U4043 ( .A(n2992),  .B(n3607),  .C(n2499), .Y(w_mem_inst_n1891));
   AOI22X1 U4044 ( .A(block[244]),  .B(n3018),  .C(w_mem_inst_w_mem[212]),  .D(n3061), .Y(n3608));
   OAI21X1 U4045 ( .A(n2992),  .B(n3609),  .C(n2446), .Y(w_mem_inst_n1890));
   AOI22X1 U4046 ( .A(block[245]),  .B(n3018),  .C(w_mem_inst_w_mem[213]),  .D(n3061), .Y(n3610));
   OAI21X1 U4047 ( .A(n2992),  .B(n3611),  .C(n2391), .Y(w_mem_inst_n1889));
   AOI22X1 U4048 ( .A(block[246]),  .B(n3018),  .C(w_mem_inst_w_mem[214]),  .D(n3061), .Y(n3612));
   OAI21X1 U4049 ( .A(n2992),  .B(n3613),  .C(n2338), .Y(w_mem_inst_n1888));
   AOI22X1 U4050 ( .A(block[247]),  .B(n3018),  .C(w_mem_inst_w_mem[215]),  .D(n3061), .Y(n3614));
   OAI21X1 U4051 ( .A(n2991),  .B(n3615),  .C(n2284), .Y(w_mem_inst_n1887));
   AOI22X1 U4052 ( .A(block[248]),  .B(n3018),  .C(w_mem_inst_w_mem[216]),  .D(n3060), .Y(n3616));
   OAI21X1 U4053 ( .A(n2991),  .B(n3617),  .C(n2241), .Y(w_mem_inst_n1886));
   AOI22X1 U4054 ( .A(block[249]),  .B(n3018),  .C(w_mem_inst_w_mem[217]),  .D(n3060), .Y(n3618));
   OAI21X1 U4055 ( .A(n2991),  .B(n3619),  .C(n2208), .Y(w_mem_inst_n1885));
   AOI22X1 U4056 ( .A(block[250]),  .B(n3018),  .C(w_mem_inst_w_mem[218]),  .D(n3060), .Y(n3620));
   OAI21X1 U4057 ( .A(n2991),  .B(n3621),  .C(n2185), .Y(w_mem_inst_n1884));
   AOI22X1 U4058 ( .A(block[251]),  .B(n3018),  .C(w_mem_inst_w_mem[219]),  .D(n3060), .Y(n3622));
   OAI21X1 U4059 ( .A(n2991),  .B(n3623),  .C(n2163), .Y(w_mem_inst_n1883));
   AOI22X1 U4060 ( .A(block[252]),  .B(n3018),  .C(w_mem_inst_w_mem[220]),  .D(n3060), .Y(n3624));
   OAI21X1 U4061 ( .A(n2991),  .B(n3625),  .C(n2324), .Y(w_mem_inst_n1882));
   AOI22X1 U4062 ( .A(block[253]),  .B(n3019),  .C(w_mem_inst_w_mem[221]),  .D(n3060), .Y(n3626));
   OAI21X1 U4063 ( .A(n2991),  .B(n3627),  .C(n2148), .Y(w_mem_inst_n1881));
   AOI22X1 U4064 ( .A(block[254]),  .B(n3019),  .C(w_mem_inst_w_mem[222]),  .D(n3060), .Y(n3628));
   OAI21X1 U4065 ( .A(n2991),  .B(n3629),  .C(n2136), .Y(w_mem_inst_n1880));
   AOI22X1 U4066 ( .A(block[255]),  .B(n3019),  .C(w_mem_inst_w_mem[223]),  .D(n3060), .Y(n3630));
   OAI21X1 U4067 ( .A(n2991),  .B(n3631),  .C(n2931), .Y(w_mem_inst_n1879));
   AOI22X1 U4068 ( .A(block[256]),  .B(n3019),  .C(w_mem_inst_w_mem[224]),  .D(n3060), .Y(n3632));
   OAI21X1 U4069 ( .A(n2991),  .B(n3633),  .C(n2873), .Y(w_mem_inst_n1878));
   AOI22X1 U4070 ( .A(block[257]),  .B(n3019),  .C(w_mem_inst_w_mem[225]),  .D(n3060), .Y(n3634));
   OAI21X1 U4071 ( .A(n2991),  .B(n3635),  .C(n2823), .Y(w_mem_inst_n1877));
   AOI22X1 U4072 ( .A(block[258]),  .B(n3019),  .C(w_mem_inst_w_mem[226]),  .D(n3060), .Y(n3636));
   OAI21X1 U4073 ( .A(n2991),  .B(n3637),  .C(n2751), .Y(w_mem_inst_n1876));
   AOI22X1 U4074 ( .A(block[259]),  .B(n3019),  .C(w_mem_inst_w_mem[227]),  .D(n3060), .Y(n3638));
   OAI21X1 U4075 ( .A(n2990),  .B(n3639),  .C(n2696), .Y(w_mem_inst_n1875));
   AOI22X1 U4076 ( .A(block[260]),  .B(n3019),  .C(w_mem_inst_w_mem[228]),  .D(n3059), .Y(n3640));
   OAI21X1 U4077 ( .A(n2990),  .B(n3641),  .C(n2627), .Y(w_mem_inst_n1874));
   AOI22X1 U4078 ( .A(block[261]),  .B(n3019),  .C(w_mem_inst_w_mem[229]),  .D(n3059), .Y(n3642));
   OAI21X1 U4079 ( .A(n2990),  .B(n3643),  .C(n2577), .Y(w_mem_inst_n1873));
   AOI22X1 U4080 ( .A(block[262]),  .B(n3019),  .C(w_mem_inst_w_mem[230]),  .D(n3059), .Y(n3644));
   OAI21X1 U4081 ( .A(n2990),  .B(n3645),  .C(n2513), .Y(w_mem_inst_n1872));
   AOI22X1 U4082 ( .A(block[263]),  .B(n3019),  .C(w_mem_inst_w_mem[231]),  .D(n3059), .Y(n3646));
   OAI21X1 U4083 ( .A(n2990),  .B(n3647),  .C(n2465), .Y(w_mem_inst_n1871));
   AOI22X1 U4084 ( .A(block[264]),  .B(n3019),  .C(w_mem_inst_w_mem[232]),  .D(n3059), .Y(n3648));
   OAI21X1 U4085 ( .A(n2990),  .B(n3649),  .C(n2407), .Y(w_mem_inst_n1870));
   AOI22X1 U4086 ( .A(block[265]),  .B(n3019),  .C(w_mem_inst_w_mem[233]),  .D(n3059), .Y(n3650));
   OAI21X1 U4087 ( .A(n2990),  .B(n3651),  .C(n2911), .Y(w_mem_inst_n1869));
   AOI22X1 U4088 ( .A(block[266]),  .B(n3020),  .C(w_mem_inst_w_mem[234]),  .D(n3059), .Y(n3652));
   OAI21X1 U4089 ( .A(n2990),  .B(n3653),  .C(n2862), .Y(w_mem_inst_n1868));
   AOI22X1 U4090 ( .A(block[267]),  .B(n3020),  .C(w_mem_inst_w_mem[235]),  .D(n3059), .Y(n3654));
   OAI21X1 U4091 ( .A(n2990),  .B(n3655),  .C(n2805), .Y(w_mem_inst_n1867));
   AOI22X1 U4092 ( .A(block[268]),  .B(n3020),  .C(w_mem_inst_w_mem[236]),  .D(n3059), .Y(n3656));
   OAI21X1 U4093 ( .A(n2990),  .B(n3657),  .C(n2740), .Y(w_mem_inst_n1866));
   AOI22X1 U4094 ( .A(block[269]),  .B(n3020),  .C(w_mem_inst_w_mem[237]),  .D(n3059), .Y(n3658));
   OAI21X1 U4095 ( .A(n2990),  .B(n3659),  .C(n2347), .Y(w_mem_inst_n1865));
   AOI22X1 U4096 ( .A(block[270]),  .B(n3020),  .C(w_mem_inst_w_mem[238]),  .D(n3059), .Y(n3660));
   OAI21X1 U4097 ( .A(n2990),  .B(n3661),  .C(n2293), .Y(w_mem_inst_n1864));
   AOI22X1 U4098 ( .A(block[271]),  .B(n3020),  .C(w_mem_inst_w_mem[239]),  .D(n3059), .Y(n3662));
   OAI21X1 U4099 ( .A(n2989),  .B(n3663),  .C(n2679), .Y(w_mem_inst_n1863));
   AOI22X1 U4100 ( .A(block[272]),  .B(n3020),  .C(w_mem_inst_w_mem[240]),  .D(n3058), .Y(n3664));
   OAI21X1 U4101 ( .A(n2989),  .B(n3665),  .C(n2617), .Y(w_mem_inst_n1862));
   AOI22X1 U4102 ( .A(block[273]),  .B(n3020),  .C(w_mem_inst_w_mem[241]),  .D(n3058), .Y(n3666));
   OAI21X1 U4103 ( .A(n2989),  .B(n3667),  .C(n2560), .Y(w_mem_inst_n1861));
   AOI22X1 U4104 ( .A(block[274]),  .B(n3020),  .C(w_mem_inst_w_mem[242]),  .D(n3058), .Y(n3668));
   OAI21X1 U4105 ( .A(n2989),  .B(n3669),  .C(n2503), .Y(w_mem_inst_n1860));
   AOI22X1 U4106 ( .A(block[275]),  .B(n3020),  .C(w_mem_inst_w_mem[243]),  .D(n3058), .Y(n3670));
   OAI21X1 U4107 ( .A(n2989),  .B(n3671),  .C(n2449), .Y(w_mem_inst_n1859));
   AOI22X1 U4108 ( .A(block[276]),  .B(n3020),  .C(w_mem_inst_w_mem[244]),  .D(n3058), .Y(n3672));
   OAI21X1 U4109 ( .A(n2989),  .B(n3673),  .C(n2394), .Y(w_mem_inst_n1858));
   AOI22X1 U4110 ( .A(block[277]),  .B(n3020),  .C(w_mem_inst_w_mem[245]),  .D(n3058), .Y(n3674));
   OAI21X1 U4111 ( .A(n2989),  .B(n3675),  .C(n2244), .Y(w_mem_inst_n1857));
   AOI22X1 U4112 ( .A(block[278]),  .B(n3020),  .C(w_mem_inst_w_mem[246]),  .D(n3058), .Y(n3676));
   OAI21X1 U4113 ( .A(n2989),  .B(n3677),  .C(n2286), .Y(w_mem_inst_n1856));
   AOI22X1 U4114 ( .A(block[279]),  .B(n3021),  .C(w_mem_inst_w_mem[247]),  .D(n3058), .Y(n3678));
   OAI21X1 U4115 ( .A(n2989),  .B(n3679),  .C(n2334), .Y(w_mem_inst_n1855));
   AOI22X1 U4116 ( .A(block[280]),  .B(n3021),  .C(w_mem_inst_w_mem[248]),  .D(n3058), .Y(n3680));
   OAI21X1 U4117 ( .A(n2989),  .B(n3681),  .C(n2211), .Y(w_mem_inst_n1854));
   AOI22X1 U4118 ( .A(block[281]),  .B(n3021),  .C(w_mem_inst_w_mem[249]),  .D(n3058), .Y(n3682));
   OAI21X1 U4119 ( .A(n2989),  .B(n3683),  .C(n2188), .Y(w_mem_inst_n1853));
   AOI22X1 U4120 ( .A(block[282]),  .B(n3021),  .C(w_mem_inst_w_mem[250]),  .D(n3058), .Y(n3684));
   OAI21X1 U4121 ( .A(n2989),  .B(n3685),  .C(n2166), .Y(w_mem_inst_n1852));
   AOI22X1 U4122 ( .A(block[283]),  .B(n3021),  .C(w_mem_inst_w_mem[251]),  .D(n3058), .Y(n3686));
   OAI21X1 U4123 ( .A(n2988),  .B(n3687),  .C(n2435), .Y(w_mem_inst_n1851));
   AOI22X1 U4124 ( .A(block[284]),  .B(n3021),  .C(w_mem_inst_w_mem[252]),  .D(n3057), .Y(n3688));
   OAI21X1 U4125 ( .A(n2988),  .B(n3689),  .C(n2379), .Y(w_mem_inst_n1850));
   AOI22X1 U4126 ( .A(block[285]),  .B(n3021),  .C(w_mem_inst_w_mem[253]),  .D(n3057), .Y(n3690));
   OAI21X1 U4127 ( .A(n2988),  .B(n3691),  .C(n2232), .Y(w_mem_inst_n1849));
   AOI22X1 U4128 ( .A(block[286]),  .B(n3021),  .C(w_mem_inst_w_mem[254]),  .D(n3057), .Y(n3692));
   OAI21X1 U4129 ( .A(n2988),  .B(n3693),  .C(n2146), .Y(w_mem_inst_n1848));
   AOI22X1 U4130 ( .A(block[287]),  .B(n3021),  .C(w_mem_inst_w_mem[255]),  .D(n3057), .Y(n3694));
   OAI21X1 U4131 ( .A(n2988),  .B(n3695),  .C(n2881), .Y(w_mem_inst_n1847));
   AOI22X1 U4132 ( .A(block[288]),  .B(n3021),  .C(w_mem_inst_w_mem[256]),  .D(n3057), .Y(n3696));
   OAI21X1 U4133 ( .A(n2988),  .B(n3697),  .C(n2923), .Y(w_mem_inst_n1846));
   AOI22X1 U4134 ( .A(block[289]),  .B(n3021),  .C(w_mem_inst_w_mem[257]),  .D(n3057), .Y(n3698));
   OAI21X1 U4135 ( .A(n2988),  .B(n3699),  .C(n2759), .Y(w_mem_inst_n1845));
   AOI22X1 U4136 ( .A(block[290]),  .B(n3021),  .C(w_mem_inst_w_mem[258]),  .D(n3057), .Y(n3700));
   OAI21X1 U4137 ( .A(n2988),  .B(n3701),  .C(n2815), .Y(w_mem_inst_n1844));
   AOI22X1 U4138 ( .A(block[291]),  .B(n3021),  .C(w_mem_inst_w_mem[259]),  .D(n3057), .Y(n3702));
   OAI21X1 U4139 ( .A(n2988),  .B(n3703),  .C(n2633), .Y(w_mem_inst_n1843));
   AOI22X1 U4140 ( .A(block[292]),  .B(n3022),  .C(w_mem_inst_w_mem[260]),  .D(n3057), .Y(n3704));
   OAI21X1 U4141 ( .A(n2988),  .B(n3705),  .C(n2689), .Y(w_mem_inst_n1842));
   AOI22X1 U4142 ( .A(block[293]),  .B(n3022),  .C(w_mem_inst_w_mem[261]),  .D(n3057), .Y(n3706));
   OAI21X1 U4143 ( .A(n2988),  .B(n3707),  .C(n2519), .Y(w_mem_inst_n1841));
   AOI22X1 U4144 ( .A(block[294]),  .B(n3022),  .C(w_mem_inst_w_mem[262]),  .D(n3057), .Y(n3708));
   OAI21X1 U4145 ( .A(n2988),  .B(n3709),  .C(n2570), .Y(w_mem_inst_n1840));
   AOI22X1 U4146 ( .A(block[295]),  .B(n3022),  .C(w_mem_inst_w_mem[263]),  .D(n3057), .Y(n3710));
   OAI21X1 U4147 ( .A(n2987),  .B(n3711),  .C(n2917), .Y(w_mem_inst_n1839));
   AOI22X1 U4148 ( .A(block[296]),  .B(n3022),  .C(w_mem_inst_w_mem[264]),  .D(n3067), .Y(n3712));
   OAI21X1 U4149 ( .A(n2987),  .B(n3713),  .C(n2868), .Y(w_mem_inst_n1838));
   AOI22X1 U4150 ( .A(block[297]),  .B(n3022),  .C(w_mem_inst_w_mem[265]),  .D(n3069), .Y(n3714));
   OAI21X1 U4151 ( .A(n2987),  .B(n3715),  .C(n2810), .Y(w_mem_inst_n1837));
   AOI22X1 U4152 ( .A(block[298]),  .B(n3022),  .C(w_mem_inst_w_mem[266]),  .D(n3068), .Y(n3716));
   OAI21X1 U4153 ( .A(n2987),  .B(n3717),  .C(n2745), .Y(w_mem_inst_n1836));
   AOI22X1 U4154 ( .A(block[299]),  .B(n3022),  .C(w_mem_inst_w_mem[267]),  .D(n3120), .Y(n3718));
   OAI21X1 U4155 ( .A(n2987),  .B(n3719),  .C(n2456), .Y(w_mem_inst_n1835));
   AOI22X1 U4156 ( .A(block[300]),  .B(n3022),  .C(w_mem_inst_w_mem[268]),  .D(n3072), .Y(n3720));
   OAI21X1 U4157 ( .A(n2987),  .B(n3721),  .C(n2401), .Y(w_mem_inst_n1834));
   AOI22X1 U4158 ( .A(block[301]),  .B(n3022),  .C(w_mem_inst_w_mem[269]),  .D(n3065), .Y(n3722));
   OAI21X1 U4159 ( .A(n2987),  .B(n3723),  .C(n2295), .Y(w_mem_inst_n1833));
   AOI22X1 U4160 ( .A(block[302]),  .B(n3022),  .C(w_mem_inst_w_mem[270]),  .D(n3063), .Y(n3724));
   OAI21X1 U4161 ( .A(n2987),  .B(n3725),  .C(n2346), .Y(w_mem_inst_n1832));
   AOI22X1 U4162 ( .A(block[303]),  .B(n3022),  .C(w_mem_inst_w_mem[271]),  .D(n3059), .Y(n3726));
   OAI21X1 U4163 ( .A(n2987),  .B(n3727),  .C(n2250), .Y(w_mem_inst_n1831));
   AOI22X1 U4164 ( .A(block[304]),  .B(n3022),  .C(w_mem_inst_w_mem[272]),  .D(n3051), .Y(n3728));
   OAI21X1 U4165 ( .A(n2987),  .B(n3729),  .C(n2673), .Y(w_mem_inst_n1830));
   AOI22X1 U4166 ( .A(block[305]),  .B(n3023),  .C(w_mem_inst_w_mem[273]),  .D(n3077), .Y(n3730));
   OAI21X1 U4167 ( .A(n2987),  .B(n3731),  .C(n2611), .Y(w_mem_inst_n1829));
   AOI22X1 U4168 ( .A(block[306]),  .B(n3023),  .C(w_mem_inst_w_mem[274]),  .D(n3052), .Y(n3732));
   OAI21X1 U4169 ( .A(n2987),  .B(n3733),  .C(n2554), .Y(w_mem_inst_n1828));
   AOI22X1 U4170 ( .A(block[307]),  .B(n3023),  .C(w_mem_inst_w_mem[275]),  .D(n3075), .Y(n3734));
   OAI21X1 U4171 ( .A(n2986),  .B(n3735),  .C(n2901), .Y(puf_8_wire_3));
   AOI22X1 U4172 ( .A(block[308]),  .B(n3023),  .C(w_mem_inst_w_mem[276]),  .D(n3056), .Y(n3736));
   OAI21X1 U4173 ( .A(n2986),  .B(n3737),  .C(n2852), .Y(w_mem_inst_n1826));
   AOI22X1 U4174 ( .A(block[309]),  .B(n3023),  .C(w_mem_inst_w_mem[277]),  .D(n3056), .Y(n3738));
   OAI21X1 U4175 ( .A(n2986),  .B(n3739),  .C(n2793), .Y(w_mem_inst_n1825));
   AOI22X1 U4176 ( .A(block[310]),  .B(n3023),  .C(w_mem_inst_w_mem[278]),  .D(n3056), .Y(n3740));
   OAI21X1 U4177 ( .A(n2986),  .B(n3741),  .C(n2729), .Y(w_mem_inst_n1824));
   AOI22X1 U4178 ( .A(block[311]),  .B(n3023),  .C(w_mem_inst_w_mem[279]),  .D(n3056), .Y(n3742));
   OAI21X1 U4179 ( .A(n2986),  .B(n3743),  .C(n2493), .Y(w_mem_inst_n1823));
   AOI22X1 U4180 ( .A(block[312]),  .B(n3023),  .C(w_mem_inst_w_mem[280]),  .D(n3056), .Y(n3744));
   OAI21X1 U4181 ( .A(n2986),  .B(n3745),  .C(n2440), .Y(w_mem_inst_n1822));
   AOI22X1 U4182 ( .A(block[313]),  .B(n3023),  .C(w_mem_inst_w_mem[281]),  .D(n3056), .Y(n3746));
   OAI21X1 U4183 ( .A(n2986),  .B(n3747),  .C(n2384), .Y(w_mem_inst_n1821));
   AOI22X1 U4184 ( .A(block[314]),  .B(n3023),  .C(w_mem_inst_w_mem[282]),  .D(n3056), .Y(n3748));
   OAI21X1 U4185 ( .A(n2986),  .B(n3749),  .C(n2328), .Y(w_mem_inst_n1820));
   AOI22X1 U4186 ( .A(block[315]),  .B(n3023),  .C(w_mem_inst_w_mem[283]),  .D(n3056), .Y(n3750));
   OAI21X1 U4187 ( .A(n2986),  .B(n3751),  .C(n2276), .Y(w_mem_inst_n1819));
   AOI22X1 U4188 ( .A(block[316]),  .B(n3023),  .C(w_mem_inst_w_mem[284]),  .D(n3056), .Y(n3752));
   OAI21X1 U4189 ( .A(n2986),  .B(n3753),  .C(n2233), .Y(w_mem_inst_n1818));
   AOI22X1 U4190 ( .A(block[317]),  .B(n3023),  .C(w_mem_inst_w_mem[285]),  .D(n3056), .Y(n3754));
   OAI21X1 U4191 ( .A(n2986),  .B(n3755),  .C(n2200), .Y(w_mem_inst_n1817));
   AOI22X1 U4192 ( .A(block[318]),  .B(n3024),  .C(w_mem_inst_w_mem[286]),  .D(n3056), .Y(n3756));
   OAI21X1 U4193 ( .A(n2986),  .B(n3757),  .C(n2177), .Y(w_mem_inst_n1816));
   AOI22X1 U4194 ( .A(block[319]),  .B(n3024),  .C(w_mem_inst_w_mem[287]),  .D(n3056), .Y(n3758));
   OAI21X1 U4195 ( .A(n2985),  .B(n3759),  .C(n2930), .Y(w_mem_inst_n1815));
   AOI22X1 U4196 ( .A(block[320]),  .B(n3024),  .C(w_mem_inst_w_mem[288]),  .D(n3055), .Y(n3760));
   OAI21X1 U4197 ( .A(n2985),  .B(n3761),  .C(n2872), .Y(w_mem_inst_n1814));
   AOI22X1 U4198 ( .A(block[321]),  .B(n3024),  .C(w_mem_inst_w_mem[289]),  .D(n3055), .Y(n3762));
   OAI21X1 U4199 ( .A(n2985),  .B(n3763),  .C(n2822), .Y(w_mem_inst_n1813));
   AOI22X1 U4200 ( .A(block[322]),  .B(n3024),  .C(w_mem_inst_w_mem[290]),  .D(n3055), .Y(n3764));
   OAI21X1 U4201 ( .A(n2985),  .B(n3765),  .C(n2700), .Y(w_mem_inst_n1812));
   AOI22X1 U4202 ( .A(block[323]),  .B(n3024),  .C(w_mem_inst_w_mem[291]),  .D(n3055), .Y(n3766));
   OAI21X1 U4203 ( .A(n2985),  .B(n3767),  .C(n2581), .Y(w_mem_inst_n1811));
   AOI22X1 U4204 ( .A(block[324]),  .B(n3024),  .C(w_mem_inst_w_mem[292]),  .D(n3055), .Y(n3768));
   OAI21X1 U4205 ( .A(n2985),  .B(n3769),  .C(n2748), .Y(w_mem_inst_n1810));
   AOI22X1 U4206 ( .A(block[325]),  .B(n3042),  .C(w_mem_inst_w_mem[293]),  .D(n3055), .Y(n3770));
   OAI21X1 U4207 ( .A(n2985),  .B(n3771),  .C(n2623), .Y(w_mem_inst_n1809));
   AOI22X1 U4208 ( .A(block[326]),  .B(n3039),  .C(w_mem_inst_w_mem[294]),  .D(n3055), .Y(n3772));
   OAI21X1 U4209 ( .A(n2985),  .B(n3773),  .C(n2512), .Y(w_mem_inst_n1808));
   AOI22X1 U4210 ( .A(block[327]),  .B(n3039),  .C(w_mem_inst_w_mem[295]),  .D(n3055), .Y(n3774));
   OAI21X1 U4211 ( .A(n2985),  .B(n3775),  .C(n2464), .Y(w_mem_inst_n1807));
   AOI22X1 U4212 ( .A(block[328]),  .B(n3039),  .C(w_mem_inst_w_mem[296]),  .D(n3055), .Y(n3776));
   OAI21X1 U4213 ( .A(n2985),  .B(n3777),  .C(n2406), .Y(w_mem_inst_n1806));
   AOI22X1 U4214 ( .A(block[329]),  .B(n3039),  .C(w_mem_inst_w_mem[297]),  .D(n3055), .Y(n3778));
   OAI21X1 U4215 ( .A(n2985),  .B(n3779),  .C(n2353), .Y(w_mem_inst_n1805));
   AOI22X1 U4216 ( .A(block[330]),  .B(n3039),  .C(w_mem_inst_w_mem[298]),  .D(n3055), .Y(n3780));
   OAI21X1 U4217 ( .A(n2985),  .B(n3781),  .C(n2300), .Y(w_mem_inst_n1804));
   AOI22X1 U4218 ( .A(block[331]),  .B(n3039),  .C(w_mem_inst_w_mem[299]),  .D(n3055), .Y(n3782));
   OAI21X1 U4219 ( .A(n2984),  .B(n3783),  .C(n2860), .Y(w_mem_inst_n1803));
   AOI22X1 U4220 ( .A(block[332]),  .B(n3039),  .C(w_mem_inst_w_mem[300]),  .D(n3054), .Y(n3784));
   OAI21X1 U4221 ( .A(n2984),  .B(n3785),  .C(n2683), .Y(w_mem_inst_n1802));
   AOI22X1 U4222 ( .A(block[333]),  .B(n3039),  .C(w_mem_inst_w_mem[301]),  .D(n3054), .Y(n3786));
   OAI21X1 U4223 ( .A(n2984),  .B(n3787),  .C(n2566), .Y(w_mem_inst_n1801));
   AOI22X1 U4224 ( .A(block[334]),  .B(n3039),  .C(w_mem_inst_w_mem[302]),  .D(n3054), .Y(n3788));
   OAI21X1 U4225 ( .A(n2984),  .B(n3789),  .C(n2252), .Y(w_mem_inst_n1800));
   AOI22X1 U4226 ( .A(block[335]),  .B(n3039),  .C(w_mem_inst_w_mem[303]),  .D(n3054), .Y(n3790));
   OAI21X1 U4227 ( .A(n2984),  .B(n3791),  .C(n2903), .Y(w_mem_inst_n1799));
   AOI22X1 U4228 ( .A(block[336]),  .B(n3040),  .C(w_mem_inst_w_mem[304]),  .D(n3054), .Y(n3792));
   OAI21X1 U4229 ( .A(n2984),  .B(n3793),  .C(n2797), .Y(w_mem_inst_n1798));
   AOI22X1 U4230 ( .A(block[337]),  .B(n3040),  .C(w_mem_inst_w_mem[305]),  .D(n3054), .Y(n3794));
   OAI21X1 U4231 ( .A(n2984),  .B(n3795),  .C(n2733), .Y(w_mem_inst_n1797));
   AOI22X1 U4232 ( .A(block[338]),  .B(n3040),  .C(w_mem_inst_w_mem[306]),  .D(n3054), .Y(n3796));
   OAI21X1 U4233 ( .A(n2984),  .B(n3797),  .C(n2608), .Y(w_mem_inst_n1796));
   AOI22X1 U4234 ( .A(block[339]),  .B(n3040),  .C(w_mem_inst_w_mem[307]),  .D(n3054), .Y(n3798));
   OAI21X1 U4235 ( .A(n2984),  .B(n3799),  .C(n2498), .Y(w_mem_inst_n1795));
   AOI22X1 U4236 ( .A(block[340]),  .B(n3040),  .C(w_mem_inst_w_mem[308]),  .D(n3054), .Y(n3800));
   OAI21X1 U4237 ( .A(n2984),  .B(n3801),  .C(n2445), .Y(w_mem_inst_n1794));
   AOI22X1 U4238 ( .A(block[341]),  .B(n3040),  .C(w_mem_inst_w_mem[309]),  .D(n3054), .Y(n3802));
   OAI21X1 U4239 ( .A(n2984),  .B(n3803),  .C(n2390), .Y(w_mem_inst_n1793));
   AOI22X1 U4240 ( .A(block[342]),  .B(n3040),  .C(w_mem_inst_w_mem[310]),  .D(n3054), .Y(n3804));
   OAI21X1 U4241 ( .A(n2984),  .B(n3805),  .C(n2337), .Y(w_mem_inst_n1792));
   AOI22X1 U4242 ( .A(block[343]),  .B(n3040),  .C(w_mem_inst_w_mem[311]),  .D(n3054), .Y(n3806));
   OAI21X1 U4243 ( .A(n2983),  .B(n3807),  .C(n2666), .Y(w_mem_inst_n1791));
   AOI22X1 U4244 ( .A(block[344]),  .B(n3040),  .C(w_mem_inst_w_mem[312]),  .D(n3071), .Y(n3808));
   OAI21X1 U4245 ( .A(n2983),  .B(n3809),  .C(n2548), .Y(w_mem_inst_n1790));
   AOI22X1 U4246 ( .A(block[345]),  .B(n3040),  .C(w_mem_inst_w_mem[313]),  .D(n3055), .Y(n3810));
   OAI21X1 U4247 ( .A(n2983),  .B(n3811),  .C(n2281), .Y(w_mem_inst_n1789));
   AOI22X1 U4248 ( .A(block[346]),  .B(n3040),  .C(w_mem_inst_w_mem[314]),  .D(n3064), .Y(n3812));
   OAI21X1 U4249 ( .A(n2983),  .B(n3813),  .C(n2237), .Y(w_mem_inst_n1788));
   AOI22X1 U4250 ( .A(block[347]),  .B(n3040),  .C(w_mem_inst_w_mem[315]),  .D(n3062), .Y(n3814));
   OAI21X1 U4251 ( .A(n2983),  .B(n3815),  .C(n2205), .Y(w_mem_inst_n1787));
   AOI22X1 U4252 ( .A(block[348]),  .B(n3040),  .C(w_mem_inst_w_mem[316]),  .D(n3057), .Y(n3816));
   OAI21X1 U4253 ( .A(n2983),  .B(n3817),  .C(n2378), .Y(w_mem_inst_n1786));
   AOI22X1 U4254 ( .A(block[349]),  .B(n3041),  .C(w_mem_inst_w_mem[317]),  .D(n3060), .Y(n3818));
   OAI21X1 U4255 ( .A(n2983),  .B(n3819),  .C(n2180), .Y(w_mem_inst_n1785));
   AOI22X1 U4256 ( .A(block[350]),  .B(n3041),  .C(w_mem_inst_w_mem[318]),  .D(n3067), .Y(n3820));
   OAI21X1 U4257 ( .A(n2983),  .B(n3821),  .C(n2158), .Y(w_mem_inst_n1784));
   AOI22X1 U4258 ( .A(block[351]),  .B(n3041),  .C(w_mem_inst_w_mem[319]),  .D(n3069), .Y(n3822));
   OAI21X1 U4259 ( .A(n2983),  .B(n3823),  .C(n2880), .Y(w_mem_inst_n1783));
   AOI22X1 U4260 ( .A(block[352]),  .B(n3041),  .C(w_mem_inst_w_mem[320]),  .D(n3068), .Y(n3824));
   OAI21X1 U4261 ( .A(n2983),  .B(n3825),  .C(n2922), .Y(w_mem_inst_n1782));
   AOI22X1 U4262 ( .A(block[353]),  .B(n3041),  .C(w_mem_inst_w_mem[321]),  .D(n3120), .Y(n3826));
   OAI21X1 U4263 ( .A(n2983),  .B(n3827),  .C(n2758), .Y(w_mem_inst_n1781));
   AOI22X1 U4264 ( .A(block[354]),  .B(n3041),  .C(w_mem_inst_w_mem[322]),  .D(n3072), .Y(n3828));
   OAI21X1 U4265 ( .A(n2983),  .B(n3829),  .C(n2814), .Y(w_mem_inst_n1780));
   AOI22X1 U4266 ( .A(block[355]),  .B(n3041),  .C(w_mem_inst_w_mem[323]),  .D(n3065), .Y(n3830));
   OAI21X1 U4267 ( .A(n2982),  .B(n3831),  .C(n2695), .Y(w_mem_inst_n1779));
   AOI22X1 U4268 ( .A(block[356]),  .B(n3041),  .C(w_mem_inst_w_mem[324]),  .D(n3053), .Y(n3832));
   OAI21X1 U4269 ( .A(n2982),  .B(n3833),  .C(n2626), .Y(w_mem_inst_n1778));
   AOI22X1 U4270 ( .A(block[357]),  .B(n3041),  .C(w_mem_inst_w_mem[325]),  .D(n3053), .Y(n3834));
   OAI21X1 U4271 ( .A(n2982),  .B(n3835),  .C(n2576), .Y(w_mem_inst_n1777));
   AOI22X1 U4272 ( .A(block[358]),  .B(n3041),  .C(w_mem_inst_w_mem[326]),  .D(n3053), .Y(n3836));
   OAI21X1 U4273 ( .A(n2982),  .B(n3837),  .C(n2469), .Y(w_mem_inst_n1776));
   AOI22X1 U4274 ( .A(block[359]),  .B(n3041),  .C(w_mem_inst_w_mem[327]),  .D(n3053), .Y(n3838));
   OAI21X1 U4275 ( .A(n2982),  .B(n3839),  .C(n2509), .Y(w_mem_inst_n1775));
   AOI22X1 U4276 ( .A(block[360]),  .B(n3041),  .C(w_mem_inst_w_mem[328]),  .D(n3053), .Y(n3840));
   OAI21X1 U4277 ( .A(n2982),  .B(n3841),  .C(n2357), .Y(w_mem_inst_n1774));
   AOI22X1 U4278 ( .A(block[361]),  .B(n3041),  .C(w_mem_inst_w_mem[329]),  .D(n3053), .Y(n3842));
   OAI21X1 U4279 ( .A(n2982),  .B(n3843),  .C(n2910), .Y(w_mem_inst_n1773));
   AOI22X1 U4280 ( .A(block[362]),  .B(n3042),  .C(w_mem_inst_w_mem[330]),  .D(n3053), .Y(n3844));
   OAI21X1 U4281 ( .A(n2982),  .B(n3845),  .C(n2861), .Y(w_mem_inst_n1772));
   AOI22X1 U4282 ( .A(block[363]),  .B(n3042),  .C(w_mem_inst_w_mem[331]),  .D(n3053), .Y(n3846));
   OAI21X1 U4283 ( .A(n2982),  .B(n3847),  .C(n2804), .Y(w_mem_inst_n1771));
   AOI22X1 U4284 ( .A(block[364]),  .B(n3042),  .C(w_mem_inst_w_mem[332]),  .D(n3053), .Y(n3848));
   OAI21X1 U4285 ( .A(n2982),  .B(n3849),  .C(n2400), .Y(w_mem_inst_n1770));
   AOI22X1 U4286 ( .A(block[365]),  .B(n3042),  .C(w_mem_inst_w_mem[333]),  .D(n3053), .Y(n3850));
   OAI21X1 U4287 ( .A(n2982),  .B(n3851),  .C(n2294), .Y(w_mem_inst_n1769));
   AOI22X1 U4288 ( .A(block[366]),  .B(n3042),  .C(w_mem_inst_w_mem[334]),  .D(n3053), .Y(n3852));
   OAI21X1 U4289 ( .A(n2982),  .B(n3853),  .C(n2213), .Y(w_mem_inst_n1768));
   AOI22X1 U4290 ( .A(block[367]),  .B(n3042),  .C(w_mem_inst_w_mem[335]),  .D(n3053), .Y(n3854));
   OAI21X1 U4291 ( .A(n2981),  .B(n3855),  .C(n2678), .Y(w_mem_inst_n1767));
   AOI22X1 U4292 ( .A(block[368]),  .B(n3042),  .C(w_mem_inst_w_mem[336]),  .D(n3057), .Y(n3856));
   OAI21X1 U4293 ( .A(n2981),  .B(n3857),  .C(n2616), .Y(w_mem_inst_n1766));
   AOI22X1 U4294 ( .A(block[369]),  .B(n3042),  .C(w_mem_inst_w_mem[337]),  .D(n3060), .Y(n3858));
   OAI21X1 U4295 ( .A(n2981),  .B(n3859),  .C(n2559), .Y(w_mem_inst_n1765));
   AOI22X1 U4296 ( .A(block[370]),  .B(n3042),  .C(w_mem_inst_w_mem[338]),  .D(n3060), .Y(n3860));
   OAI21X1 U4297 ( .A(n2981),  .B(n3861),  .C(n2502), .Y(w_mem_inst_n1764));
   AOI22X1 U4298 ( .A(block[371]),  .B(n3042),  .C(w_mem_inst_w_mem[339]),  .D(n3067), .Y(n3862));
   OAI21X1 U4299 ( .A(n2981),  .B(n3863),  .C(n2448), .Y(w_mem_inst_n1763));
   AOI22X1 U4300 ( .A(block[372]),  .B(n3042),  .C(w_mem_inst_w_mem[340]),  .D(n3069), .Y(n3864));
   OAI21X1 U4301 ( .A(n2981),  .B(n3865),  .C(n2341), .Y(w_mem_inst_n1762));
   AOI22X1 U4302 ( .A(block[373]),  .B(n3042),  .C(w_mem_inst_w_mem[341]),  .D(n3068), .Y(n3866));
   OAI21X1 U4303 ( .A(n2981),  .B(n3867),  .C(n2730), .Y(w_mem_inst_n1761));
   AOI22X1 U4304 ( .A(block[374]),  .B(n3020),  .C(w_mem_inst_w_mem[342]),  .D(n3120), .Y(n3868));
   OAI21X1 U4305 ( .A(n2981),  .B(n3869),  .C(n2388), .Y(w_mem_inst_n1760));
   AOI22X1 U4306 ( .A(block[375]),  .B(n3030),  .C(w_mem_inst_w_mem[343]),  .D(n3072), .Y(n3870));
   OAI21X1 U4307 ( .A(n2981),  .B(n3871),  .C(n2283), .Y(w_mem_inst_n1759));
   AOI22X1 U4308 ( .A(block[376]),  .B(n3028),  .C(w_mem_inst_w_mem[344]),  .D(n3065), .Y(n3872));
   OAI21X1 U4309 ( .A(n2981),  .B(n3873),  .C(n2240), .Y(w_mem_inst_n1758));
   AOI22X1 U4310 ( .A(block[377]),  .B(n3024),  .C(w_mem_inst_w_mem[345]),  .D(n3063), .Y(n3874));
   OAI21X1 U4311 ( .A(n2981),  .B(n3875),  .C(n2207), .Y(w_mem_inst_n1757));
   AOI22X1 U4312 ( .A(block[378]),  .B(n3013),  .C(w_mem_inst_w_mem[346]),  .D(n3059), .Y(n3876));
   OAI21X1 U4313 ( .A(n2981),  .B(n3877),  .C(n2184), .Y(w_mem_inst_n1756));
   AOI22X1 U4314 ( .A(block[379]),  .B(n3021),  .C(w_mem_inst_w_mem[347]),  .D(n3051), .Y(n3878));
   OAI21X1 U4315 ( .A(n2999),  .B(n3879),  .C(n2434), .Y(w_mem_inst_n1755));
   AOI22X1 U4316 ( .A(block[380]),  .B(n3022),  .C(w_mem_inst_w_mem[348]),  .D(n3052), .Y(n3880));
   OAI21X1 U4317 ( .A(n3005),  .B(n3881),  .C(n2323), .Y(w_mem_inst_n1754));
   AOI22X1 U4318 ( .A(block[381]),  .B(n3035),  .C(w_mem_inst_w_mem[349]),  .D(n3052), .Y(n3882));
   OAI21X1 U4319 ( .A(n2981),  .B(n3883),  .C(n2160), .Y(w_mem_inst_n1753));
   AOI22X1 U4320 ( .A(block[382]),  .B(n3040),  .C(w_mem_inst_w_mem[350]),  .D(n3052), .Y(n3884));
   OAI21X1 U4321 ( .A(n3003),  .B(n3885),  .C(n2145), .Y(w_mem_inst_n1752));
   AOI22X1 U4322 ( .A(block[383]),  .B(n3025),  .C(w_mem_inst_w_mem[351]),  .D(n3052), .Y(n3886));
   OAI21X1 U4323 ( .A(n2993),  .B(n3887),  .C(n2929), .Y(w_mem_inst_n1751));
   AOI22X1 U4324 ( .A(block[384]),  .B(n3031),  .C(w_mem_inst_w_mem[352]),  .D(n3052), .Y(n3888));
   OAI21X1 U4325 ( .A(n2992),  .B(n3889),  .C(n2871), .Y(w_mem_inst_n1750));
   AOI22X1 U4326 ( .A(block[385]),  .B(n3042),  .C(w_mem_inst_w_mem[353]),  .D(n3052), .Y(n3890));
   OAI21X1 U4327 ( .A(n3009),  .B(n3891),  .C(n2821), .Y(w_mem_inst_n1749));
   AOI22X1 U4328 ( .A(block[386]),  .B(n3017),  .C(w_mem_inst_w_mem[354]),  .D(n3052), .Y(n3892));
   OAI21X1 U4329 ( .A(n2998),  .B(n3893),  .C(n2750), .Y(w_mem_inst_n1748));
   AOI22X1 U4330 ( .A(block[387]),  .B(n3015),  .C(w_mem_inst_w_mem[355]),  .D(n3052), .Y(n3894));
   OAI21X1 U4331 ( .A(n2987),  .B(n3895),  .C(n2632), .Y(w_mem_inst_n1747));
   AOI22X1 U4332 ( .A(block[388]),  .B(n3016),  .C(w_mem_inst_w_mem[356]),  .D(n3052), .Y(n3896));
   OAI21X1 U4333 ( .A(n2994),  .B(n3897),  .C(n2688), .Y(w_mem_inst_n1746));
   AOI22X1 U4334 ( .A(block[389]),  .B(n3032),  .C(w_mem_inst_w_mem[357]),  .D(n3052), .Y(n3898));
   OAI21X1 U4335 ( .A(n2989),  .B(n3899),  .C(n2518), .Y(w_mem_inst_n1745));
   AOI22X1 U4336 ( .A(block[390]),  .B(n3036),  .C(w_mem_inst_w_mem[358]),  .D(n3052), .Y(n3900));
   OAI21X1 U4337 ( .A(n2985),  .B(n3901),  .C(n2569), .Y(w_mem_inst_n1744));
   AOI22X1 U4338 ( .A(block[391]),  .B(n3019),  .C(w_mem_inst_w_mem[359]),  .D(n3052), .Y(n3902));
   OAI21X1 U4339 ( .A(n3001),  .B(n3903),  .C(n2916), .Y(w_mem_inst_n1743));
   AOI22X1 U4340 ( .A(block[392]),  .B(n3026),  .C(w_mem_inst_w_mem[360]),  .D(n3076), .Y(n3904));
   OAI21X1 U4341 ( .A(n3002),  .B(n3905),  .C(n2867), .Y(w_mem_inst_n1742));
   AOI22X1 U4342 ( .A(block[393]),  .B(n3014),  .C(w_mem_inst_w_mem[361]),  .D(n3053), .Y(n3906));
   OAI21X1 U4343 ( .A(n2986),  .B(n3907),  .C(n2809), .Y(w_mem_inst_n1741));
   AOI22X1 U4344 ( .A(block[394]),  .B(n3020),  .C(w_mem_inst_w_mem[362]),  .D(n3071), .Y(n3908));
   OAI21X1 U4345 ( .A(n3011),  .B(n3909),  .C(n2457), .Y(w_mem_inst_n1740));
   AOI22X1 U4346 ( .A(block[395]),  .B(n3030),  .C(w_mem_inst_w_mem[363]),  .D(n3055), .Y(n3910));
   OAI21X1 U4347 ( .A(n2990),  .B(n3911),  .C(n2402), .Y(w_mem_inst_n1739));
   AOI22X1 U4348 ( .A(block[396]),  .B(n3028),  .C(w_mem_inst_w_mem[364]),  .D(n3064), .Y(n3912));
   OAI21X1 U4349 ( .A(n3008),  .B(n3913),  .C(n2349), .Y(w_mem_inst_n1738));
   AOI22X1 U4350 ( .A(block[397]),  .B(n3024),  .C(w_mem_inst_w_mem[365]),  .D(n3062), .Y(n3914));
   OAI21X1 U4351 ( .A(n2983),  .B(n3915),  .C(n2256), .Y(w_mem_inst_n1737));
   AOI22X1 U4352 ( .A(block[398]),  .B(n3013),  .C(w_mem_inst_w_mem[366]),  .D(n3057), .Y(n3916));
   OAI21X1 U4353 ( .A(n3000),  .B(n3917),  .C(n2292), .Y(w_mem_inst_n1736));
   AOI22X1 U4354 ( .A(block[399]),  .B(n3021),  .C(w_mem_inst_w_mem[367]),  .D(n3060), .Y(n3918));
   OAI21X1 U4355 ( .A(n2991),  .B(n3919),  .C(n2734), .Y(w_mem_inst_n1735));
   AOI22X1 U4356 ( .A(block[400]),  .B(n3040),  .C(w_mem_inst_w_mem[368]),  .D(n3067), .Y(n3920));
   OAI21X1 U4357 ( .A(n3006),  .B(n3921),  .C(n2672), .Y(w_mem_inst_n1734));
   AOI22X1 U4358 ( .A(block[401]),  .B(n3025),  .C(w_mem_inst_w_mem[369]),  .D(n3069), .Y(n3922));
   OAI21X1 U4359 ( .A(n2984),  .B(n3923),  .C(n2610), .Y(w_mem_inst_n1733));
   AOI22X1 U4360 ( .A(block[402]),  .B(n3031),  .C(w_mem_inst_w_mem[370]),  .D(n3068), .Y(n3924));
   OAI21X1 U4361 ( .A(n2982),  .B(n3925),  .C(n2553), .Y(w_mem_inst_n1732));
   AOI22X1 U4362 ( .A(block[403]),  .B(n3042),  .C(w_mem_inst_w_mem[371]),  .D(n3120), .Y(n3926));
   OAI21X1 U4363 ( .A(n3001),  .B(n3927),  .C(n2900), .Y(w_mem_inst_n1731));
   AOI22X1 U4364 ( .A(block[404]),  .B(n3017),  .C(w_mem_inst_w_mem[372]),  .D(n3056), .Y(n3928));
   OAI21X1 U4365 ( .A(n3002),  .B(n3929),  .C(n2851), .Y(w_mem_inst_n1730));
   AOI22X1 U4366 ( .A(block[405]),  .B(n3033),  .C(w_mem_inst_w_mem[373]),  .D(n3074), .Y(n3930));
   OAI21X1 U4367 ( .A(n2986),  .B(n3931),  .C(n2792), .Y(w_mem_inst_n1729));
   AOI22X1 U4368 ( .A(block[406]),  .B(n3023),  .C(w_mem_inst_w_mem[374]),  .D(n3056), .Y(n3932));
   OAI21X1 U4369 ( .A(n3011),  .B(n3933),  .C(n2494), .Y(w_mem_inst_n1728));
   AOI22X1 U4370 ( .A(block[407]),  .B(n3036),  .C(w_mem_inst_w_mem[375]),  .D(n3078), .Y(n3934));
   OAI21X1 U4371 ( .A(n2990),  .B(n3935),  .C(n2441), .Y(w_mem_inst_n1727));
   AOI22X1 U4372 ( .A(block[408]),  .B(n3029),  .C(w_mem_inst_w_mem[376]),  .D(n3076), .Y(n3936));
   OAI21X1 U4373 ( .A(n3008),  .B(n3937),  .C(n2385), .Y(w_mem_inst_n1726));
   AOI22X1 U4374 ( .A(block[409]),  .B(n3027),  .C(w_mem_inst_w_mem[377]),  .D(n3053), .Y(n3938));
   OAI21X1 U4375 ( .A(n2983),  .B(n3939),  .C(n2330), .Y(w_mem_inst_n1725));
   AOI22X1 U4376 ( .A(block[410]),  .B(n3038),  .C(w_mem_inst_w_mem[378]),  .D(n3071), .Y(n3940));
   OAI21X1 U4377 ( .A(n3000),  .B(n3941),  .C(n2278), .Y(w_mem_inst_n1724));
   AOI22X1 U4378 ( .A(block[411]),  .B(n3034),  .C(w_mem_inst_w_mem[379]),  .D(n3055), .Y(n3942));
   OAI21X1 U4379 ( .A(n2991),  .B(n3943),  .C(n2234), .Y(w_mem_inst_n1723));
   AOI22X1 U4380 ( .A(block[412]),  .B(n3018),  .C(w_mem_inst_w_mem[380]),  .D(n3064), .Y(n3944));
   OAI21X1 U4381 ( .A(n3006),  .B(n3945),  .C(n2727), .Y(w_mem_inst_n1722));
   AOI22X1 U4382 ( .A(block[413]),  .B(n3050),  .C(w_mem_inst_w_mem[381]),  .D(n3062), .Y(n3946));
   OAI21X1 U4383 ( .A(n2984),  .B(n3947),  .C(n2664), .Y(w_mem_inst_n1721));
   AOI22X1 U4384 ( .A(block[414]),  .B(n3050),  .C(w_mem_inst_w_mem[382]),  .D(n3076), .Y(n3948));
   OAI21X1 U4385 ( .A(n2982),  .B(n3949),  .C(n2602), .Y(w_mem_inst_n1720));
   AOI22X1 U4386 ( .A(block[415]),  .B(n3050),  .C(w_mem_inst_w_mem[383]),  .D(n3057), .Y(n3950));
   OAI21X1 U4387 ( .A(n3003),  .B(n3951),  .C(n2879), .Y(w_mem_inst_n1719));
   AOI22X1 U4388 ( .A(block[416]),  .B(n3050),  .C(w_mem_inst_w_mem[384]),  .D(n3051), .Y(n3952));
   OAI21X1 U4389 ( .A(n2997),  .B(n3953),  .C(n2921), .Y(w_mem_inst_n1718));
   AOI22X1 U4390 ( .A(block[417]),  .B(n3050),  .C(w_mem_inst_w_mem[385]),  .D(n3077), .Y(n3954));
   OAI21X1 U4391 ( .A(n2993),  .B(n3955),  .C(n2757), .Y(w_mem_inst_n1717));
   AOI22X1 U4392 ( .A(block[418]),  .B(n3039),  .C(w_mem_inst_w_mem[386]),  .D(n3052), .Y(n3956));
   OAI21X1 U4393 ( .A(n2992),  .B(n3957),  .C(n2813), .Y(w_mem_inst_n1716));
   AOI22X1 U4394 ( .A(block[419]),  .B(n3039),  .C(w_mem_inst_w_mem[387]),  .D(n3075), .Y(n3958));
   OAI21X1 U4395 ( .A(n3009),  .B(n3959),  .C(n2694), .Y(w_mem_inst_n1715));
   AOI22X1 U4396 ( .A(block[420]),  .B(n3038),  .C(w_mem_inst_w_mem[388]),  .D(n3070), .Y(n3960));
   OAI21X1 U4397 ( .A(n2998),  .B(n3961),  .C(n2625), .Y(w_mem_inst_n1714));
   AOI22X1 U4398 ( .A(block[421]),  .B(n3038),  .C(w_mem_inst_w_mem[389]),  .D(n3058), .Y(n3962));
   OAI21X1 U4399 ( .A(n2987),  .B(n3963),  .C(n2575), .Y(w_mem_inst_n1713));
   AOI22X1 U4400 ( .A(block[422]),  .B(n3038),  .C(w_mem_inst_w_mem[390]),  .D(n3066), .Y(n3964));
   OAI21X1 U4401 ( .A(n2994),  .B(n3965),  .C(n2511), .Y(w_mem_inst_n1712));
   AOI22X1 U4402 ( .A(block[423]),  .B(n3038),  .C(w_mem_inst_w_mem[391]),  .D(n3054), .Y(n3966));
   OAI21X1 U4403 ( .A(n2989),  .B(n3967),  .C(n2463), .Y(w_mem_inst_n1711));
   AOI22X1 U4404 ( .A(block[424]),  .B(n3038),  .C(w_mem_inst_w_mem[392]),  .D(n3061), .Y(n3968));
   OAI21X1 U4405 ( .A(n2985),  .B(n3969),  .C(n2405), .Y(w_mem_inst_n1710));
   AOI22X1 U4406 ( .A(block[425]),  .B(n3038),  .C(w_mem_inst_w_mem[393]),  .D(n3073), .Y(n3970));
   OAI21X1 U4407 ( .A(n2996),  .B(n3971),  .C(n2352), .Y(w_mem_inst_n1709));
   AOI22X1 U4408 ( .A(block[426]),  .B(n3038),  .C(w_mem_inst_w_mem[394]),  .D(n3080), .Y(n3972));
   OAI21X1 U4409 ( .A(n2996),  .B(n3973),  .C(n2299), .Y(w_mem_inst_n1708));
   AOI22X1 U4410 ( .A(block[427]),  .B(n3038),  .C(w_mem_inst_w_mem[395]),  .D(n3079), .Y(n3974));
   OAI21X1 U4411 ( .A(n2990),  .B(n3975),  .C(n2905), .Y(w_mem_inst_n1707));
   AOI22X1 U4412 ( .A(block[428]),  .B(n3038),  .C(w_mem_inst_w_mem[396]),  .D(n3066), .Y(n3976));
   OAI21X1 U4413 ( .A(n3008),  .B(n3977),  .C(n2855), .Y(w_mem_inst_n1706));
   AOI22X1 U4414 ( .A(block[429]),  .B(n3038),  .C(w_mem_inst_w_mem[397]),  .D(n3054), .Y(n3978));
   OAI21X1 U4415 ( .A(n2983),  .B(n3979),  .C(n2800), .Y(w_mem_inst_n1705));
   AOI22X1 U4416 ( .A(block[430]),  .B(n3038),  .C(w_mem_inst_w_mem[398]),  .D(n3061), .Y(n3980));
   OAI21X1 U4417 ( .A(n3000),  .B(n3981),  .C(n2735), .Y(w_mem_inst_n1704));
   AOI22X1 U4418 ( .A(block[431]),  .B(n3038),  .C(w_mem_inst_w_mem[399]),  .D(n3073), .Y(n3982));
   OAI21X1 U4419 ( .A(n2991),  .B(n3983),  .C(n2249), .Y(w_mem_inst_n1703));
   AOI22X1 U4420 ( .A(block[432]),  .B(n3038),  .C(w_mem_inst_w_mem[400]),  .D(n3063), .Y(n3984));
   OAI21X1 U4421 ( .A(n3006),  .B(n3985),  .C(n2615), .Y(w_mem_inst_n1702));
   AOI22X1 U4422 ( .A(block[433]),  .B(n3037),  .C(w_mem_inst_w_mem[401]),  .D(n3065), .Y(n3986));
   OAI21X1 U4423 ( .A(n2984),  .B(n3987),  .C(n2671), .Y(w_mem_inst_n1701));
   AOI22X1 U4424 ( .A(block[434]),  .B(n3037),  .C(w_mem_inst_w_mem[402]),  .D(n3080), .Y(n3988));
   OAI21X1 U4425 ( .A(n2982),  .B(n3989),  .C(n2501), .Y(w_mem_inst_n1700));
   AOI22X1 U4426 ( .A(block[435]),  .B(n3037),  .C(w_mem_inst_w_mem[403]),  .D(n3079), .Y(n3990));
   OAI21X1 U4427 ( .A(n2997),  .B(n3991),  .C(n2552), .Y(puf_9_wire_3));
   AOI22X1 U4428 ( .A(block[436]),  .B(n3037),  .C(w_mem_inst_w_mem[404]),  .D(n3074), .Y(n3992));
   OAI21X1 U4429 ( .A(n3010),  .B(n3993),  .C(n2444), .Y(w_mem_inst_n1698));
   AOI22X1 U4430 ( .A(block[437]),  .B(n3037),  .C(w_mem_inst_w_mem[405]),  .D(n3074), .Y(n3994));
   OAI21X1 U4431 ( .A(n3007),  .B(n3995),  .C(n2389), .Y(w_mem_inst_n1697));
   AOI22X1 U4432 ( .A(block[438]),  .B(n3037),  .C(w_mem_inst_w_mem[406]),  .D(n3056), .Y(n3996));
   OAI21X1 U4433 ( .A(n2999),  .B(n3997),  .C(n2336), .Y(w_mem_inst_n1696));
   AOI22X1 U4434 ( .A(block[439]),  .B(n3037),  .C(w_mem_inst_w_mem[407]),  .D(n3078), .Y(n3998));
   OAI21X1 U4435 ( .A(n2994),  .B(n3999),  .C(n2282), .Y(w_mem_inst_n1695));
   AOI22X1 U4436 ( .A(block[440]),  .B(n3037),  .C(w_mem_inst_w_mem[408]),  .D(n3051), .Y(n4000));
   OAI21X1 U4437 ( .A(n2989),  .B(n4001),  .C(n2239), .Y(w_mem_inst_n1694));
   AOI22X1 U4438 ( .A(block[441]),  .B(n3037),  .C(w_mem_inst_w_mem[409]),  .D(n3051), .Y(n4002));
   OAI21X1 U4439 ( .A(n2986),  .B(n4003),  .C(n2206), .Y(w_mem_inst_n1693));
   AOI22X1 U4440 ( .A(block[442]),  .B(n3037),  .C(w_mem_inst_w_mem[410]),  .D(n3051), .Y(n4004));
   OAI21X1 U4441 ( .A(n2985),  .B(n4005),  .C(n2183), .Y(w_mem_inst_n1692));
   AOI22X1 U4442 ( .A(block[443]),  .B(n3037),  .C(w_mem_inst_w_mem[411]),  .D(n3051), .Y(n4006));
   OAI21X1 U4443 ( .A(n2996),  .B(n4007),  .C(n2162), .Y(w_mem_inst_n1691));
   AOI22X1 U4444 ( .A(block[444]),  .B(n3037),  .C(w_mem_inst_w_mem[412]),  .D(n3051), .Y(n4008));
   OAI21X1 U4445 ( .A(n3004),  .B(n4009),  .C(n2150), .Y(w_mem_inst_n1690));
   AOI22X1 U4446 ( .A(block[445]),  .B(n3037),  .C(w_mem_inst_w_mem[413]),  .D(n3051), .Y(n4010));
   OAI21X1 U4447 ( .A(n3004),  .B(n4011),  .C(n2322), .Y(w_mem_inst_n1689));
   AOI22X1 U4448 ( .A(block[446]),  .B(n3032),  .C(w_mem_inst_w_mem[414]),  .D(n3051), .Y(n4012));
   OAI21X1 U4449 ( .A(n2988),  .B(n4013),  .C(n2135), .Y(w_mem_inst_n1688));
   AOI22X1 U4450 ( .A(block[447]),  .B(n3039),  .C(w_mem_inst_w_mem[415]),  .D(n3051), .Y(n4014));
   OAI21X1 U4451 ( .A(n2995),  .B(n4015),  .C(n2928), .Y(w_mem_inst_n1687));
   AOI22X1 U4452 ( .A(block[448]),  .B(n3016),  .C(w_mem_inst_w_mem[416]),  .D(n3051), .Y(n4016));
   OAI21X1 U4453 ( .A(n3001),  .B(n4017),  .C(n2870), .Y(w_mem_inst_n1686));
   AOI22X1 U4454 ( .A(block[449]),  .B(n3015),  .C(w_mem_inst_w_mem[417]),  .D(n3051), .Y(n4018));
   OAI21X1 U4455 ( .A(n3002),  .B(n4019),  .C(n2820), .Y(w_mem_inst_n1685));
   AOI22X1 U4456 ( .A(block[450]),  .B(n3046),  .C(w_mem_inst_w_mem[418]),  .D(n3051), .Y(n4020));
   OAI21X1 U4457 ( .A(n3004),  .B(n4021),  .C(n2749), .Y(w_mem_inst_n1684));
   AOI22X1 U4458 ( .A(block[451]),  .B(n3046),  .C(w_mem_inst_w_mem[419]),  .D(n3051), .Y(n4022));
   OAI21X1 U4459 ( .A(n3010),  .B(n4023),  .C(n2631), .Y(w_mem_inst_n1683));
   AOI22X1 U4460 ( .A(block[452]),  .B(n3044),  .C(w_mem_inst_w_mem[420]),  .D(n3052), .Y(n4024));
   OAI21X1 U4461 ( .A(n3007),  .B(n4025),  .C(n2687), .Y(w_mem_inst_n1682));
   AOI22X1 U4462 ( .A(block[453]),  .B(n3047),  .C(w_mem_inst_w_mem[421]),  .D(n3075), .Y(n4026));
   OAI21X1 U4463 ( .A(n2999),  .B(n4027),  .C(n2517), .Y(w_mem_inst_n1681));
   AOI22X1 U4464 ( .A(block[454]),  .B(n3045),  .C(w_mem_inst_w_mem[422]),  .D(n3070), .Y(n4028));
   OAI21X1 U4465 ( .A(n3005),  .B(n4029),  .C(n2568), .Y(w_mem_inst_n1680));
   AOI22X1 U4466 ( .A(block[455]),  .B(n3043),  .C(w_mem_inst_w_mem[423]),  .D(n3058), .Y(n4030));
   OAI21X1 U4467 ( .A(n2981),  .B(n4031),  .C(n2411), .Y(w_mem_inst_n1679));
   AOI22X1 U4468 ( .A(block[456]),  .B(n3050),  .C(w_mem_inst_w_mem[424]),  .D(n3066), .Y(n4032));
   OAI21X1 U4469 ( .A(n3003),  .B(n4033),  .C(n2460), .Y(w_mem_inst_n1678));
   AOI22X1 U4470 ( .A(block[457]),  .B(n3041),  .C(w_mem_inst_w_mem[425]),  .D(n3054), .Y(n4034));
   OAI21X1 U4471 ( .A(n3010),  .B(n4035),  .C(n2304), .Y(w_mem_inst_n1677));
   AOI22X1 U4472 ( .A(block[458]),  .B(n3048),  .C(w_mem_inst_w_mem[426]),  .D(n3061), .Y(n4036));
   OAI21X1 U4473 ( .A(n2993),  .B(n4037),  .C(n2909), .Y(w_mem_inst_n1676));
   AOI22X1 U4474 ( .A(block[459]),  .B(n3040),  .C(w_mem_inst_w_mem[427]),  .D(n3073), .Y(n4038));
   OAI21X1 U4475 ( .A(n3005),  .B(n4039),  .C(n2859), .Y(w_mem_inst_n1675));
   AOI22X1 U4476 ( .A(block[460]),  .B(n3035),  .C(w_mem_inst_w_mem[428]),  .D(n3059), .Y(n4040));
   OAI21X1 U4477 ( .A(n2992),  .B(n4041),  .C(n2803), .Y(w_mem_inst_n1674));
   AOI22X1 U4478 ( .A(block[461]),  .B(n3022),  .C(w_mem_inst_w_mem[429]),  .D(n3063), .Y(n4042));
   OAI21X1 U4479 ( .A(n3009),  .B(n4043),  .C(n2738), .Y(w_mem_inst_n1673));
   AOI22X1 U4480 ( .A(block[462]),  .B(n3021),  .C(w_mem_inst_w_mem[430]),  .D(n3070), .Y(n4044));
   OAI21X1 U4481 ( .A(n2998),  .B(n4045),  .C(n2345), .Y(w_mem_inst_n1672));
   AOI22X1 U4482 ( .A(block[463]),  .B(n3013),  .C(w_mem_inst_w_mem[431]),  .D(n3080), .Y(n4046));
   OAI21X1 U4483 ( .A(n2981),  .B(n4047),  .C(n2677), .Y(w_mem_inst_n1671));
   AOI22X1 U4484 ( .A(block[464]),  .B(n3024),  .C(w_mem_inst_w_mem[432]),  .D(n3078), .Y(n4048));
   OAI21X1 U4485 ( .A(n3003),  .B(n4049),  .C(n2563), .Y(w_mem_inst_n1670));
   AOI22X1 U4486 ( .A(block[465]),  .B(n3035),  .C(w_mem_inst_w_mem[433]),  .D(n3074), .Y(n4050));
   OAI21X1 U4487 ( .A(n2989),  .B(n4051),  .C(n2609), .Y(w_mem_inst_n1669));
   AOI22X1 U4488 ( .A(block[466]),  .B(n3028),  .C(w_mem_inst_w_mem[434]),  .D(n3056), .Y(n4052));
   OAI21X1 U4489 ( .A(n3011),  .B(n4053),  .C(n2453), .Y(w_mem_inst_n1668));
   AOI22X1 U4490 ( .A(block[467]),  .B(n3030),  .C(w_mem_inst_w_mem[435]),  .D(n3078), .Y(n4054));
   OAI21X1 U4491 ( .A(n2985),  .B(n4055),  .C(n2497), .Y(w_mem_inst_n1667));
   AOI22X1 U4492 ( .A(block[468]),  .B(n3020),  .C(w_mem_inst_w_mem[436]),  .D(n3076), .Y(n4056));
   OAI21X1 U4493 ( .A(n2997),  .B(n4057),  .C(n2393), .Y(w_mem_inst_n1666));
   AOI22X1 U4494 ( .A(block[469]),  .B(n3014),  .C(w_mem_inst_w_mem[437]),  .D(n3053), .Y(n4058));
   OAI21X1 U4495 ( .A(n2987),  .B(n4059),  .C(n2288), .Y(w_mem_inst_n1665));
   AOI22X1 U4496 ( .A(block[470]),  .B(n3026),  .C(w_mem_inst_w_mem[438]),  .D(n3079), .Y(n4060));
   OAI21X1 U4497 ( .A(n2996),  .B(n4061),  .C(n2243), .Y(w_mem_inst_n1664));
   AOI22X1 U4498 ( .A(block[471]),  .B(n3019),  .C(w_mem_inst_w_mem[439]),  .D(n3071), .Y(n4062));
   OAI21X1 U4499 ( .A(n2988),  .B(n4063),  .C(n2333), .Y(w_mem_inst_n1663));
   AOI22X1 U4500 ( .A(block[472]),  .B(n3026),  .C(w_mem_inst_w_mem[440]),  .D(n3055), .Y(n4064));
   OAI21X1 U4501 ( .A(n3004),  .B(n4065),  .C(n2210), .Y(w_mem_inst_n1662));
   AOI22X1 U4502 ( .A(block[473]),  .B(n3019),  .C(w_mem_inst_w_mem[441]),  .D(n3064), .Y(n4066));
   OAI21X1 U4503 ( .A(n2988),  .B(n4067),  .C(n2187), .Y(w_mem_inst_n1661));
   AOI22X1 U4504 ( .A(block[474]),  .B(n3033),  .C(w_mem_inst_w_mem[442]),  .D(n3062), .Y(n4068));
   OAI21X1 U4505 ( .A(n2995),  .B(n4069),  .C(n2165), .Y(w_mem_inst_n1660));
   AOI22X1 U4506 ( .A(block[475]),  .B(n3032),  .C(w_mem_inst_w_mem[443]),  .D(n3053), .Y(n4070));
   OAI21X1 U4507 ( .A(n3002),  .B(n4071),  .C(n2433), .Y(w_mem_inst_n1659));
   AOI22X1 U4508 ( .A(block[476]),  .B(n3023),  .C(w_mem_inst_w_mem[444]),  .D(n3077), .Y(n4072));
   OAI21X1 U4509 ( .A(n2988),  .B(n4073),  .C(n2377), .Y(w_mem_inst_n1658));
   AOI22X1 U4510 ( .A(block[477]),  .B(n3037),  .C(w_mem_inst_w_mem[445]),  .D(n3052), .Y(n4074));
   OAI21X1 U4511 ( .A(n2986),  .B(n4075),  .C(n2272), .Y(w_mem_inst_n1657));
   AOI22X1 U4512 ( .A(block[478]),  .B(n3016),  .C(w_mem_inst_w_mem[446]),  .D(n3075), .Y(n4076));
   OAI21X1 U4513 ( .A(n3011),  .B(n4077),  .C(n2229), .Y(w_mem_inst_n1656));
   AOI22X1 U4514 ( .A(block[479]),  .B(n3015),  .C(w_mem_inst_w_mem[447]),  .D(n3070), .Y(n4078));
   OAI21X1 U4515 ( .A(n2990),  .B(n4079),  .C(n2878), .Y(w_mem_inst_n1655));
   AOI22X1 U4516 ( .A(block[480]),  .B(n3044),  .C(w_mem_inst_w_mem[448]),  .D(n3058), .Y(n4080));
   OAI21X1 U4517 ( .A(n3008),  .B(n4081),  .C(n2920), .Y(w_mem_inst_n1654));
   AOI22X1 U4518 ( .A(block[481]),  .B(n3044),  .C(w_mem_inst_w_mem[449]),  .D(n3066), .Y(n4082));
   OAI21X1 U4519 ( .A(n2983),  .B(n4083),  .C(n2756), .Y(w_mem_inst_n1653));
   AOI22X1 U4520 ( .A(block[482]),  .B(n3047),  .C(w_mem_inst_w_mem[450]),  .D(n3054), .Y(n4084));
   OAI21X1 U4521 ( .A(n3000),  .B(n4085),  .C(n2812), .Y(w_mem_inst_n1652));
   AOI22X1 U4522 ( .A(block[483]),  .B(n3045),  .C(w_mem_inst_w_mem[451]),  .D(n3061), .Y(n4086));
   OAI21X1 U4523 ( .A(n2991),  .B(n4087),  .C(n2693), .Y(w_mem_inst_n1651));
   AOI22X1 U4524 ( .A(block[484]),  .B(n3043),  .C(w_mem_inst_w_mem[452]),  .D(n3073), .Y(n4088));
   OAI21X1 U4525 ( .A(n3006),  .B(n4089),  .C(n2624), .Y(w_mem_inst_n1650));
   AOI22X1 U4526 ( .A(block[485]),  .B(n3025),  .C(w_mem_inst_w_mem[453]),  .D(n3072), .Y(n4090));
   OAI21X1 U4527 ( .A(n2984),  .B(n4091),  .C(n2574), .Y(w_mem_inst_n1649));
   AOI22X1 U4528 ( .A(block[486]),  .B(n3040),  .C(w_mem_inst_w_mem[454]),  .D(n3080), .Y(n4092));
   OAI21X1 U4529 ( .A(n2982),  .B(n4093),  .C(n2510), .Y(w_mem_inst_n1648));
   AOI22X1 U4530 ( .A(block[487]),  .B(n3035),  .C(w_mem_inst_w_mem[455]),  .D(n3079), .Y(n4094));
   OAI21X1 U4531 ( .A(n2983),  .B(n4095),  .C(n2915), .Y(w_mem_inst_n1647));
   AOI22X1 U4532 ( .A(block[488]),  .B(n3022),  .C(w_mem_inst_w_mem[456]),  .D(n3070), .Y(n4096));
   OAI21X1 U4533 ( .A(n3000),  .B(n4097),  .C(n2866), .Y(w_mem_inst_n1646));
   AOI22X1 U4534 ( .A(block[489]),  .B(n3021),  .C(w_mem_inst_w_mem[457]),  .D(n3058), .Y(n4098));
   OAI21X1 U4535 ( .A(n2991),  .B(n4099),  .C(n2808), .Y(w_mem_inst_n1645));
   AOI22X1 U4536 ( .A(block[490]),  .B(n3013),  .C(w_mem_inst_w_mem[458]),  .D(n3066), .Y(n4100));
   OAI21X1 U4537 ( .A(n3006),  .B(n4101),  .C(n2744), .Y(w_mem_inst_n1644));
   AOI22X1 U4538 ( .A(block[491]),  .B(n3025),  .C(w_mem_inst_w_mem[459]),  .D(n3054), .Y(n4102));
   OAI21X1 U4539 ( .A(n2984),  .B(n4103),  .C(n2685), .Y(w_mem_inst_n1643));
   AOI22X1 U4540 ( .A(block[492]),  .B(n3024),  .C(w_mem_inst_w_mem[460]),  .D(n3061), .Y(n4104));
   OAI21X1 U4541 ( .A(n2982),  .B(n4105),  .C(n2455), .Y(w_mem_inst_n1642));
   AOI22X1 U4542 ( .A(block[493]),  .B(n3022),  .C(w_mem_inst_w_mem[461]),  .D(n3073), .Y(n4106));
   OAI21X1 U4543 ( .A(n3001),  .B(n4107),  .C(n2399), .Y(w_mem_inst_n1641));
   AOI22X1 U4544 ( .A(block[494]),  .B(n3028),  .C(w_mem_inst_w_mem[462]),  .D(n3051), .Y(n4108));
   OAI21X1 U4545 ( .A(n2997),  .B(n4109),  .C(n2291), .Y(w_mem_inst_n1640));
   AOI22X1 U4546 ( .A(block[495]),  .B(n3030),  .C(w_mem_inst_w_mem[463]),  .D(n3059), .Y(n4110));
   OAI21X1 U4547 ( .A(n3010),  .B(n4111),  .C(n2344), .Y(w_mem_inst_n1639));
   AOI22X1 U4548 ( .A(block[496]),  .B(n3020),  .C(w_mem_inst_w_mem[464]),  .D(n3058), .Y(n4112));
   OAI21X1 U4549 ( .A(n3007),  .B(n4113),  .C(n2248), .Y(w_mem_inst_n1638));
   AOI22X1 U4550 ( .A(block[497]),  .B(n3014),  .C(w_mem_inst_w_mem[465]),  .D(n3080), .Y(n4114));
   OAI21X1 U4551 ( .A(n2999),  .B(n4115),  .C(n2558), .Y(w_mem_inst_n1637));
   AOI22X1 U4552 ( .A(block[498]),  .B(n3039),  .C(w_mem_inst_w_mem[466]),  .D(n3079), .Y(n4116));
   OAI21X1 U4553 ( .A(n3005),  .B(n4117),  .C(n2607), .Y(w_mem_inst_n1636));
   AOI22X1 U4554 ( .A(block[499]),  .B(n3037),  .C(w_mem_inst_w_mem[467]),  .D(n3077), .Y(n4118));
   OAI21X1 U4555 ( .A(n2996),  .B(n4119),  .C(n2899), .Y(w_mem_inst_n1635));
   AOI22X1 U4556 ( .A(block[500]),  .B(n3018),  .C(w_mem_inst_w_mem[468]),  .D(n3120), .Y(n4120));
   OAI21X1 U4557 ( .A(n2995),  .B(n4121),  .C(n2850), .Y(w_mem_inst_n1634));
   AOI22X1 U4558 ( .A(block[501]),  .B(n3034),  .C(w_mem_inst_w_mem[469]),  .D(n3120), .Y(n4122));
   OAI21X1 U4559 ( .A(n3004),  .B(n4123),  .C(n2791), .Y(w_mem_inst_n1633));
   AOI22X1 U4560 ( .A(block[502]),  .B(n3038),  .C(w_mem_inst_w_mem[470]),  .D(n3120), .Y(n4124));
   OAI21X1 U4561 ( .A(n2988),  .B(n4125),  .C(n2728), .Y(w_mem_inst_n1632));
   AOI22X1 U4562 ( .A(block[503]),  .B(n3027),  .C(w_mem_inst_w_mem[471]),  .D(n3120), .Y(n4126));
   OAI21X1 U4563 ( .A(n2995),  .B(n4127),  .C(n2665), .Y(w_mem_inst_n1631));
   AOI22X1 U4564 ( .A(block[504]),  .B(n3029),  .C(w_mem_inst_w_mem[472]),  .D(n3072), .Y(n4128));
   OAI21X1 U4565 ( .A(n3001),  .B(n4129),  .C(n2492), .Y(w_mem_inst_n1630));
   AOI22X1 U4566 ( .A(block[505]),  .B(n3036),  .C(w_mem_inst_w_mem[473]),  .D(n3065), .Y(n4130));
   OAI21X1 U4567 ( .A(n3002),  .B(n4131),  .C(n2439), .Y(w_mem_inst_n1629));
   AOI22X1 U4568 ( .A(block[506]),  .B(n3023),  .C(w_mem_inst_w_mem[474]),  .D(n3063), .Y(n4132));
   OAI21X1 U4569 ( .A(n2995),  .B(n4133),  .C(n2383), .Y(w_mem_inst_n1628));
   AOI22X1 U4570 ( .A(block[507]),  .B(n3033),  .C(w_mem_inst_w_mem[475]),  .D(n3059), .Y(n4134));
   OAI21X1 U4571 ( .A(n2986),  .B(n4135),  .C(n2327), .Y(w_mem_inst_n1627));
   AOI22X1 U4572 ( .A(block[508]),  .B(n3017),  .C(w_mem_inst_w_mem[476]),  .D(n3051), .Y(n4136));
   OAI21X1 U4573 ( .A(n3011),  .B(n4137),  .C(n2274), .Y(w_mem_inst_n1626));
   AOI22X1 U4574 ( .A(block[509]),  .B(n3042),  .C(w_mem_inst_w_mem[477]),  .D(n3077), .Y(n4138));
   OAI21X1 U4575 ( .A(n2990),  .B(n4139),  .C(n2231), .Y(w_mem_inst_n1625));
   AOI22X1 U4576 ( .A(block[510]),  .B(n3031),  .C(w_mem_inst_w_mem[478]),  .D(n3052), .Y(n4140));
   OAI21X1 U4577 ( .A(n3008),  .B(n4141),  .C(n2199), .Y(w_mem_inst_n1624));
   AOI22X1 U4578 ( .A(block[511]),  .B(n3036),  .C(w_mem_inst_w_mem[479]),  .D(n3075), .Y(n4142));
   INVX1 U4579 ( .A(n4143), .Y(n3120));
   NAND3X1 U4580 ( .A(n3116),  .B(n3100),  .C(n2957), .Y(n4143));
   NAND3X1 U4581 ( .A(n3116),  .B(n3100),  .C(n4144), .Y(n3117));
   FAX1 U4582 ( .A(n3221),  .B(n3217),  .C(w_mem_inst_w_mem[42]), .YS(w_mem_inst_N639));
   FAX1 U4583 ( .A(n3223),  .B(n3219),  .C(w_mem_inst_w_mem[43]), .YS(w_mem_inst_N638));
   FAX1 U4584 ( .A(n3225),  .B(n3221),  .C(w_mem_inst_w_mem[44]), .YS(w_mem_inst_N637));
   FAX1 U4585 ( .A(n3227),  .B(n3223),  .C(w_mem_inst_w_mem[45]), .YS(w_mem_inst_N636));
   FAX1 U4586 ( .A(n3229),  .B(n3225),  .C(w_mem_inst_w_mem[46]), .YS(w_mem_inst_N635));
   FAX1 U4587 ( .A(n3231),  .B(n3227),  .C(w_mem_inst_w_mem[47]), .YS(w_mem_inst_N634));
   FAX1 U4588 ( .A(n3233),  .B(n3229),  .C(w_mem_inst_w_mem[48]), .YS(w_mem_inst_N633));
   FAX1 U4589 ( .A(n3235),  .B(n3231),  .C(w_mem_inst_w_mem[49]), .YS(w_mem_inst_N632));
   FAX1 U4590 ( .A(n3237),  .B(n3233),  .C(w_mem_inst_w_mem[50]), .YS(w_mem_inst_N631));
   FAX1 U4591 ( .A(n3239),  .B(n3235),  .C(w_mem_inst_w_mem[51]), .YS(w_mem_inst_N630));
   FAX1 U4592 ( .A(n3241),  .B(n3237),  .C(w_mem_inst_w_mem[52]), .YS(w_mem_inst_N629));
   FAX1 U4593 ( .A(n3243),  .B(n3239),  .C(w_mem_inst_w_mem[53]), .YS(w_mem_inst_N628));
   FAX1 U4594 ( .A(n3245),  .B(n3241),  .C(w_mem_inst_w_mem[54]), .YS(w_mem_inst_N627));
   FAX1 U4595 ( .A(n3243),  .B(n3229),  .C(w_mem_inst_w_mem[32]), .YS(w_mem_inst_N626));
   FAX1 U4596 ( .A(n3245),  .B(n3231),  .C(w_mem_inst_w_mem[33]), .YS(w_mem_inst_N625));
   FAX1 U4597 ( .A(n3187),  .B(n3233),  .C(w_mem_inst_w_mem[32]), .YS(w_mem_inst_N624));
   FAX1 U4598 ( .A(n3189),  .B(n3235),  .C(w_mem_inst_w_mem[33]), .YS(w_mem_inst_N623));
   FAX1 U4599 ( .A(n3191),  .B(n3187),  .C(w_mem_inst_w_mem[59]), .YS(w_mem_inst_N622));
   FAX1 U4600 ( .A(n3193),  .B(n3189),  .C(w_mem_inst_w_mem[60]), .YS(w_mem_inst_N621));
   FAX1 U4601 ( .A(n3195),  .B(n3191),  .C(w_mem_inst_w_mem[61]), .YS(w_mem_inst_N620));
   FAX1 U4602 ( .A(n3197),  .B(n3193),  .C(w_mem_inst_w_mem[62]), .YS(w_mem_inst_N619));
   FAX1 U4603 ( .A(n3199),  .B(n3195),  .C(w_mem_inst_w_mem[63]), .YS(w_mem_inst_N618));
   XNOR2X1 U4604 ( .A(n3201),  .B(w_mem_inst_w_mem[39]), .Y(w_mem_inst_N617));
   XNOR2X1 U4605 ( .A(n3199),  .B(w_mem_inst_w_mem[42]), .Y(w_mem_inst_N616));
   XNOR2X1 U4606 ( .A(n3201),  .B(w_mem_inst_w_mem[43]), .Y(w_mem_inst_N615));
   XNOR2X1 U4607 ( .A(n3207),  .B(w_mem_inst_w_mem[42]), .Y(w_mem_inst_N614));
   XNOR2X1 U4608 ( .A(n3209),  .B(w_mem_inst_w_mem[43]), .Y(w_mem_inst_N613));
   XNOR2X1 U4609 ( .A(n3211),  .B(w_mem_inst_w_mem[44]), .Y(w_mem_inst_N612));
   XNOR2X1 U4610 ( .A(n3213),  .B(w_mem_inst_w_mem[45]), .Y(w_mem_inst_N611));
   XNOR2X1 U4611 ( .A(n3215),  .B(w_mem_inst_w_mem[46]), .Y(w_mem_inst_N610));
   XNOR2X1 U4612 ( .A(n3217),  .B(w_mem_inst_w_mem[47]), .Y(w_mem_inst_N609));
   XNOR2X1 U4613 ( .A(n3219),  .B(w_mem_inst_w_mem[48]), .Y(w_mem_inst_N608));
   FAX1 U4614 ( .A(n4029),  .B(n4021),  .C(w_mem_inst_w_mem[466]), .YS(w_mem_inst_N607));
   FAX1 U4615 ( .A(n4031),  .B(n4023),  .C(w_mem_inst_w_mem[467]), .YS(w_mem_inst_N606));
   FAX1 U4616 ( .A(n4033),  .B(n4025),  .C(w_mem_inst_w_mem[468]), .YS(w_mem_inst_N605));
   FAX1 U4617 ( .A(n4027),  .B(n4057),  .C(w_mem_inst_w_mem[458]), .YS(w_mem_inst_N604));
   FAX1 U4618 ( .A(n4029),  .B(n4059),  .C(w_mem_inst_w_mem[459]), .YS(w_mem_inst_N603));
   FAX1 U4619 ( .A(n4031),  .B(n4061),  .C(w_mem_inst_w_mem[460]), .YS(w_mem_inst_N602));
   FAX1 U4620 ( .A(n4033),  .B(n4063),  .C(w_mem_inst_w_mem[461]), .YS(w_mem_inst_N601));
   FAX1 U4621 ( .A(n4065),  .B(n4043),  .C(w_mem_inst_w_mem[458]), .YS(w_mem_inst_N600));
   FAX1 U4622 ( .A(n4067),  .B(n4045),  .C(w_mem_inst_w_mem[459]), .YS(w_mem_inst_N599));
   FAX1 U4623 ( .A(n4069),  .B(n4047),  .C(w_mem_inst_w_mem[460]), .YS(w_mem_inst_N598));
   FAX1 U4624 ( .A(n4071),  .B(n4049),  .C(w_mem_inst_w_mem[461]), .YS(w_mem_inst_N597));
   FAX1 U4625 ( .A(n4073),  .B(n4051),  .C(w_mem_inst_w_mem[462]), .YS(w_mem_inst_N596));
   FAX1 U4626 ( .A(n4075),  .B(n4053),  .C(w_mem_inst_w_mem[463]), .YS(w_mem_inst_N595));
   FAX1 U4627 ( .A(n4077),  .B(n4055),  .C(w_mem_inst_w_mem[464]), .YS(w_mem_inst_N594));
   FAX1 U4628 ( .A(n4057),  .B(n4049),  .C(w_mem_inst_w_mem[448]), .YS(w_mem_inst_N593));
   FAX1 U4629 ( .A(n4059),  .B(n4017),  .C(w_mem_inst_w_mem[466]), .YS(w_mem_inst_N592));
   FAX1 U4630 ( .A(n4019),  .B(n4061),  .C(w_mem_inst_w_mem[467]), .YS(w_mem_inst_N591));
   FAX1 U4631 ( .A(n4021),  .B(n4063),  .C(w_mem_inst_w_mem[468]), .YS(w_mem_inst_N590));
   FAX1 U4632 ( .A(n4023),  .B(n4065),  .C(w_mem_inst_w_mem[469]), .YS(w_mem_inst_N589));
   FAX1 U4633 ( .A(n4025),  .B(n4067),  .C(w_mem_inst_w_mem[470]), .YS(w_mem_inst_N588));
   FAX1 U4634 ( .A(n4027),  .B(n4069),  .C(w_mem_inst_w_mem[471]), .YS(w_mem_inst_N587));
   FAX1 U4635 ( .A(n4029),  .B(n4071),  .C(w_mem_inst_w_mem[472]), .YS(w_mem_inst_N586));
   FAX1 U4636 ( .A(n4031),  .B(n4073),  .C(w_mem_inst_w_mem[473]), .YS(w_mem_inst_N585));
   FAX1 U4637 ( .A(n4033),  .B(n4075),  .C(w_mem_inst_w_mem[474]), .YS(w_mem_inst_N584));
   FAX1 U4638 ( .A(n4077),  .B(n4069),  .C(w_mem_inst_w_mem[458]), .YS(w_mem_inst_N583));
   FAX1 U4639 ( .A(n4071),  .B(n4037),  .C(w_mem_inst_w_mem[448]), .YS(w_mem_inst_N582));
   FAX1 U4640 ( .A(n4073),  .B(n4017),  .C(w_mem_inst_w_mem[460]), .YS(w_mem_inst_N581));
   FAX1 U4641 ( .A(n4075),  .B(n4019),  .C(w_mem_inst_w_mem[461]), .YS(w_mem_inst_N580));
   FAX1 U4642 ( .A(n4021),  .B(n4077),  .C(w_mem_inst_w_mem[462]), .YS(w_mem_inst_N579));
   XNOR2X1 U4643 ( .A(n4023),  .B(w_mem_inst_w_mem[463]), .Y(w_mem_inst_N578));
   XNOR2X1 U4644 ( .A(n4025),  .B(w_mem_inst_w_mem[464]), .Y(w_mem_inst_N577));
   XNOR2X1 U4645 ( .A(n4027),  .B(w_mem_inst_w_mem[465]), .Y(w_mem_inst_N576));
   NAND3X1 U4646 ( .A(n4149),  .B(n4150),  .C(n4151), .Y(n4148));
   AOI22X1 U4647 ( .A(n2121),  .B(n3841),  .C(n2125),  .D(n3969), .Y(n4151));
   INVX1 U4648 ( .A(w_mem_inst_w_mem[425]), .Y(n3969));
   INVX1 U4649 ( .A(w_mem_inst_w_mem[361]), .Y(n3841));
   NAND2X1 U4650 ( .A(n2119),  .B(n4097), .Y(n4150));
   INVX1 U4651 ( .A(w_mem_inst_w_mem[489]), .Y(n4097));
   NAND3X1 U4652 ( .A(n4155),  .B(n4156),  .C(n4157), .Y(n4147));
   AOI22X1 U4653 ( .A(n4158),  .B(n4033),  .C(n2123),  .D(n3713), .Y(n4157));
   INVX1 U4654 ( .A(w_mem_inst_w_mem[297]), .Y(n3713));
   INVX1 U4655 ( .A(w_mem_inst_w_mem[457]), .Y(n4033));
   NAND2X1 U4656 ( .A(n3106),  .B(n3649), .Y(n4156));
   INVX1 U4657 ( .A(w_mem_inst_w_mem[265]), .Y(n3649));
   AOI22X1 U4658 ( .A(n4160),  .B(n3777),  .C(n4161),  .D(n3905), .Y(n4155));
   INVX1 U4659 ( .A(w_mem_inst_w_mem[393]), .Y(n3905));
   INVX1 U4660 ( .A(w_mem_inst_w_mem[329]), .Y(n3777));
   NAND3X1 U4661 ( .A(n4162),  .B(n4163),  .C(n4164), .Y(n4145));
   AND2X1 U4662 ( .A(n4165),  .B(n4166), .Y(n4164));
   AOI22X1 U4663 ( .A(n4158),  .B(n3521),  .C(n2123),  .D(n3201), .Y(n4166));
   INVX1 U4664 ( .A(w_mem_inst_w_mem[41]), .Y(n3201));
   INVX1 U4665 ( .A(w_mem_inst_w_mem[201]), .Y(n3521));
   AOI22X1 U4666 ( .A(n2121),  .B(n3329),  .C(n2125),  .D(n3457), .Y(n4165));
   INVX1 U4667 ( .A(w_mem_inst_w_mem[169]), .Y(n3457));
   INVX1 U4668 ( .A(w_mem_inst_w_mem[105]), .Y(n3329));
   OAI21X1 U4669 ( .A(n4160),  .B(n3393),  .C(n4167), .Y(n4163));
   AOI21X1 U4670 ( .A(w_mem_inst_w_mem[73]),  .B(n2958),  .C(n4169), .Y(n4167));
   INVX1 U4671 ( .A(w_mem_inst_w_mem[137]), .Y(n3393));
   AOI22X1 U4672 ( .A(n2119),  .B(n3585),  .C(n2117),  .D(n4171), .Y(n4162));
   NAND2X1 U4673 ( .A(n4442),  .B(w_mem_inst_w_mem[9]), .Y(n4171));
   INVX1 U4674 ( .A(w_mem_inst_w_mem[233]), .Y(n3585));
   NAND3X1 U4675 ( .A(n4149),  .B(n4176),  .C(n4177), .Y(n4175));
   AOI22X1 U4676 ( .A(n2121),  .B(n3839),  .C(n2125),  .D(n3967), .Y(n4177));
   INVX1 U4677 ( .A(w_mem_inst_w_mem[424]), .Y(n3967));
   INVX1 U4678 ( .A(w_mem_inst_w_mem[360]), .Y(n3839));
   NAND2X1 U4679 ( .A(n2119),  .B(n4095), .Y(n4176));
   INVX1 U4680 ( .A(w_mem_inst_w_mem[488]), .Y(n4095));
   NAND3X1 U4681 ( .A(n4178),  .B(n4179),  .C(n4180), .Y(n4174));
   AOI22X1 U4682 ( .A(n4158),  .B(n4031),  .C(n2123),  .D(n3711), .Y(n4180));
   INVX1 U4683 ( .A(w_mem_inst_w_mem[296]), .Y(n3711));
   INVX1 U4684 ( .A(w_mem_inst_w_mem[456]), .Y(n4031));
   NAND2X1 U4685 ( .A(n3106),  .B(n3647), .Y(n4179));
   INVX1 U4686 ( .A(w_mem_inst_w_mem[264]), .Y(n3647));
   AOI22X1 U4687 ( .A(n4160),  .B(n3775),  .C(n4161),  .D(n3903), .Y(n4178));
   INVX1 U4688 ( .A(w_mem_inst_w_mem[392]), .Y(n3903));
   INVX1 U4689 ( .A(w_mem_inst_w_mem[328]), .Y(n3775));
   NAND3X1 U4690 ( .A(n4181),  .B(n4182),  .C(n4183), .Y(n4172));
   AND2X1 U4691 ( .A(n4184),  .B(n4185), .Y(n4183));
   AOI22X1 U4692 ( .A(n4158),  .B(n3519),  .C(n2123),  .D(n3199), .Y(n4185));
   INVX1 U4693 ( .A(w_mem_inst_w_mem[40]), .Y(n3199));
   INVX1 U4694 ( .A(w_mem_inst_w_mem[200]), .Y(n3519));
   AOI22X1 U4695 ( .A(n2121),  .B(n3327),  .C(n2125),  .D(n3455), .Y(n4184));
   INVX1 U4696 ( .A(w_mem_inst_w_mem[168]), .Y(n3455));
   INVX1 U4697 ( .A(w_mem_inst_w_mem[104]), .Y(n3327));
   OAI21X1 U4698 ( .A(n4160),  .B(n3391),  .C(n4186), .Y(n4182));
   AOI21X1 U4699 ( .A(w_mem_inst_w_mem[72]),  .B(n2958),  .C(n4169), .Y(n4186));
   INVX1 U4700 ( .A(w_mem_inst_w_mem[136]), .Y(n3391));
   AOI22X1 U4701 ( .A(n2119),  .B(n3583),  .C(n2117),  .D(n4187), .Y(n4181));
   NAND2X1 U4702 ( .A(n4442),  .B(w_mem_inst_w_mem[8]), .Y(n4187));
   INVX1 U4703 ( .A(w_mem_inst_w_mem[232]), .Y(n3583));
   NAND3X1 U4704 ( .A(n4149),  .B(n4192),  .C(n4193), .Y(n4191));
   AOI22X1 U4705 ( .A(n2121),  .B(n3837),  .C(n2125),  .D(n3965), .Y(n4193));
   INVX1 U4706 ( .A(w_mem_inst_w_mem[423]), .Y(n3965));
   INVX1 U4707 ( .A(w_mem_inst_w_mem[359]), .Y(n3837));
   NAND2X1 U4708 ( .A(n2119),  .B(n4093), .Y(n4192));
   INVX1 U4709 ( .A(w_mem_inst_w_mem[487]), .Y(n4093));
   NAND3X1 U4710 ( .A(n4194),  .B(n4195),  .C(n4196), .Y(n4190));
   AOI22X1 U4711 ( .A(n4158),  .B(n4029),  .C(n2123),  .D(n3709), .Y(n4196));
   INVX1 U4712 ( .A(w_mem_inst_w_mem[295]), .Y(n3709));
   INVX1 U4713 ( .A(w_mem_inst_w_mem[455]), .Y(n4029));
   NAND2X1 U4714 ( .A(n3106),  .B(n3645), .Y(n4195));
   INVX1 U4715 ( .A(w_mem_inst_w_mem[263]), .Y(n3645));
   AOI22X1 U4716 ( .A(n4160),  .B(n3773),  .C(n4161),  .D(n3901), .Y(n4194));
   INVX1 U4717 ( .A(w_mem_inst_w_mem[391]), .Y(n3901));
   INVX1 U4718 ( .A(w_mem_inst_w_mem[327]), .Y(n3773));
   NAND3X1 U4719 ( .A(n4197),  .B(n4198),  .C(n4199), .Y(n4188));
   AND2X1 U4720 ( .A(n4200),  .B(n4201), .Y(n4199));
   AOI22X1 U4721 ( .A(n4158),  .B(n3517),  .C(n2123),  .D(n3197), .Y(n4201));
   INVX1 U4722 ( .A(w_mem_inst_w_mem[39]), .Y(n3197));
   INVX1 U4723 ( .A(w_mem_inst_w_mem[199]), .Y(n3517));
   AOI22X1 U4724 ( .A(n2121),  .B(n3325),  .C(n2125),  .D(n3453), .Y(n4200));
   INVX1 U4725 ( .A(w_mem_inst_w_mem[167]), .Y(n3453));
   INVX1 U4726 ( .A(w_mem_inst_w_mem[103]), .Y(n3325));
   OAI21X1 U4727 ( .A(n4160),  .B(n3389),  .C(n4202), .Y(n4198));
   AOI21X1 U4728 ( .A(w_mem_inst_w_mem[71]),  .B(n2958),  .C(n4169), .Y(n4202));
   INVX1 U4729 ( .A(w_mem_inst_w_mem[135]), .Y(n3389));
   AOI22X1 U4730 ( .A(n2119),  .B(n3581),  .C(n2117),  .D(n4203), .Y(n4197));
   NAND2X1 U4731 ( .A(n4442),  .B(w_mem_inst_w_mem[7]), .Y(n4203));
   INVX1 U4732 ( .A(w_mem_inst_w_mem[231]), .Y(n3581));
   NAND3X1 U4733 ( .A(n4149),  .B(n4208),  .C(n4209), .Y(n4207));
   AOI22X1 U4734 ( .A(n2121),  .B(n3835),  .C(n2125),  .D(n3963), .Y(n4209));
   INVX1 U4735 ( .A(w_mem_inst_w_mem[422]), .Y(n3963));
   INVX1 U4736 ( .A(w_mem_inst_w_mem[358]), .Y(n3835));
   NAND2X1 U4737 ( .A(n2119),  .B(n4091), .Y(n4208));
   INVX1 U4738 ( .A(w_mem_inst_w_mem[486]), .Y(n4091));
   NAND3X1 U4739 ( .A(n4210),  .B(n4211),  .C(n4212), .Y(n4206));
   AOI22X1 U4740 ( .A(n4158),  .B(n4027),  .C(n2123),  .D(n3707), .Y(n4212));
   INVX1 U4741 ( .A(w_mem_inst_w_mem[294]), .Y(n3707));
   INVX1 U4742 ( .A(w_mem_inst_w_mem[454]), .Y(n4027));
   NAND2X1 U4743 ( .A(n3106),  .B(n3643), .Y(n4211));
   INVX1 U4744 ( .A(w_mem_inst_w_mem[262]), .Y(n3643));
   AOI22X1 U4745 ( .A(n4160),  .B(n3771),  .C(n4161),  .D(n3899), .Y(n4210));
   INVX1 U4746 ( .A(w_mem_inst_w_mem[390]), .Y(n3899));
   INVX1 U4747 ( .A(w_mem_inst_w_mem[326]), .Y(n3771));
   NAND3X1 U4748 ( .A(n4213),  .B(n4214),  .C(n4215), .Y(n4204));
   AND2X1 U4749 ( .A(n4216),  .B(n4217), .Y(n4215));
   AOI22X1 U4750 ( .A(n4158),  .B(n3515),  .C(n2123),  .D(n3195), .Y(n4217));
   INVX1 U4751 ( .A(w_mem_inst_w_mem[38]), .Y(n3195));
   INVX1 U4752 ( .A(w_mem_inst_w_mem[198]), .Y(n3515));
   AOI22X1 U4753 ( .A(n2121),  .B(n3323),  .C(n2125),  .D(n3451), .Y(n4216));
   INVX1 U4754 ( .A(w_mem_inst_w_mem[166]), .Y(n3451));
   INVX1 U4755 ( .A(w_mem_inst_w_mem[102]), .Y(n3323));
   OAI21X1 U4756 ( .A(n4160),  .B(n3387),  .C(n4218), .Y(n4214));
   AOI21X1 U4757 ( .A(w_mem_inst_w_mem[70]),  .B(n2958),  .C(n4169), .Y(n4218));
   INVX1 U4758 ( .A(w_mem_inst_w_mem[134]), .Y(n3387));
   AOI22X1 U4759 ( .A(n2119),  .B(n3579),  .C(n2117),  .D(n4219), .Y(n4213));
   NAND2X1 U4760 ( .A(n4442),  .B(w_mem_inst_w_mem[6]), .Y(n4219));
   INVX1 U4761 ( .A(w_mem_inst_w_mem[230]), .Y(n3579));
   NAND3X1 U4762 ( .A(n4149),  .B(n4224),  .C(n4225), .Y(n4223));
   AOI22X1 U4763 ( .A(n2121),  .B(n3833),  .C(n2125),  .D(n3961), .Y(n4225));
   INVX1 U4764 ( .A(w_mem_inst_w_mem[421]), .Y(n3961));
   INVX1 U4765 ( .A(w_mem_inst_w_mem[357]), .Y(n3833));
   NAND2X1 U4766 ( .A(n2119),  .B(n4089), .Y(n4224));
   INVX1 U4767 ( .A(w_mem_inst_w_mem[485]), .Y(n4089));
   NAND3X1 U4768 ( .A(n4226),  .B(n4227),  .C(n4228), .Y(n4222));
   AOI22X1 U4769 ( .A(n4158),  .B(n4025),  .C(n2123),  .D(n3705), .Y(n4228));
   INVX1 U4770 ( .A(w_mem_inst_w_mem[293]), .Y(n3705));
   INVX1 U4771 ( .A(w_mem_inst_w_mem[453]), .Y(n4025));
   NAND2X1 U4772 ( .A(n3106),  .B(n3641), .Y(n4227));
   INVX1 U4773 ( .A(w_mem_inst_w_mem[261]), .Y(n3641));
   AOI22X1 U4774 ( .A(n4160),  .B(n3769),  .C(n4161),  .D(n3897), .Y(n4226));
   INVX1 U4775 ( .A(w_mem_inst_w_mem[389]), .Y(n3897));
   INVX1 U4776 ( .A(w_mem_inst_w_mem[325]), .Y(n3769));
   NAND3X1 U4777 ( .A(n4229),  .B(n4230),  .C(n4231), .Y(n4220));
   AND2X1 U4778 ( .A(n4232),  .B(n4233), .Y(n4231));
   AOI22X1 U4779 ( .A(n4158),  .B(n3513),  .C(n2123),  .D(n3193), .Y(n4233));
   INVX1 U4780 ( .A(w_mem_inst_w_mem[37]), .Y(n3193));
   INVX1 U4781 ( .A(w_mem_inst_w_mem[197]), .Y(n3513));
   AOI22X1 U4782 ( .A(n2121),  .B(n3321),  .C(n2125),  .D(n3449), .Y(n4232));
   INVX1 U4783 ( .A(w_mem_inst_w_mem[165]), .Y(n3449));
   INVX1 U4784 ( .A(w_mem_inst_w_mem[101]), .Y(n3321));
   OAI21X1 U4785 ( .A(n4160),  .B(n3385),  .C(n4234), .Y(n4230));
   AOI21X1 U4786 ( .A(w_mem_inst_w_mem[69]),  .B(n2958),  .C(n4169), .Y(n4234));
   INVX1 U4787 ( .A(w_mem_inst_w_mem[133]), .Y(n3385));
   AOI22X1 U4788 ( .A(n2119),  .B(n3577),  .C(n2117),  .D(n4235), .Y(n4229));
   NAND2X1 U4789 ( .A(n4442),  .B(w_mem_inst_w_mem[5]), .Y(n4235));
   INVX1 U4790 ( .A(w_mem_inst_w_mem[229]), .Y(n3577));
   NAND3X1 U4791 ( .A(n4149),  .B(n4240),  .C(n4241), .Y(n4239));
   AOI22X1 U4792 ( .A(n2121),  .B(n3831),  .C(n2125),  .D(n3959), .Y(n4241));
   INVX1 U4793 ( .A(w_mem_inst_w_mem[420]), .Y(n3959));
   INVX1 U4794 ( .A(w_mem_inst_w_mem[356]), .Y(n3831));
   NAND2X1 U4795 ( .A(n2119),  .B(n4087), .Y(n4240));
   INVX1 U4796 ( .A(w_mem_inst_w_mem[484]), .Y(n4087));
   NAND3X1 U4797 ( .A(n4242),  .B(n4243),  .C(n4244), .Y(n4238));
   AOI22X1 U4798 ( .A(n4158),  .B(n4023),  .C(n2123),  .D(n3703), .Y(n4244));
   INVX1 U4799 ( .A(w_mem_inst_w_mem[292]), .Y(n3703));
   INVX1 U4800 ( .A(w_mem_inst_w_mem[452]), .Y(n4023));
   NAND2X1 U4801 ( .A(n3106),  .B(n3639), .Y(n4243));
   INVX1 U4802 ( .A(w_mem_inst_w_mem[260]), .Y(n3639));
   AOI22X1 U4803 ( .A(n4160),  .B(n3767),  .C(n4161),  .D(n3895), .Y(n4242));
   INVX1 U4804 ( .A(w_mem_inst_w_mem[388]), .Y(n3895));
   INVX1 U4805 ( .A(w_mem_inst_w_mem[324]), .Y(n3767));
   NAND3X1 U4806 ( .A(n4245),  .B(n4246),  .C(n4247), .Y(n4236));
   AND2X1 U4807 ( .A(n4248),  .B(n4249), .Y(n4247));
   AOI22X1 U4808 ( .A(n4158),  .B(n3511),  .C(n2123),  .D(n3191), .Y(n4249));
   INVX1 U4809 ( .A(w_mem_inst_w_mem[36]), .Y(n3191));
   INVX1 U4810 ( .A(w_mem_inst_w_mem[196]), .Y(n3511));
   AOI22X1 U4811 ( .A(n2121),  .B(n3319),  .C(n2125),  .D(n3447), .Y(n4248));
   INVX1 U4812 ( .A(w_mem_inst_w_mem[164]), .Y(n3447));
   INVX1 U4813 ( .A(w_mem_inst_w_mem[100]), .Y(n3319));
   OAI21X1 U4814 ( .A(n4160),  .B(n3383),  .C(n4250), .Y(n4246));
   AOI21X1 U4815 ( .A(w_mem_inst_w_mem[68]),  .B(n2958),  .C(n4169), .Y(n4250));
   INVX1 U4816 ( .A(w_mem_inst_w_mem[132]), .Y(n3383));
   AOI22X1 U4817 ( .A(n2119),  .B(n3575),  .C(n2117),  .D(n4251), .Y(n4245));
   NAND2X1 U4818 ( .A(n4442),  .B(w_mem_inst_w_mem[4]), .Y(n4251));
   INVX1 U4819 ( .A(w_mem_inst_w_mem[228]), .Y(n3575));
   NAND3X1 U4820 ( .A(n4149),  .B(n4256),  .C(n4257), .Y(n4255));
   AOI22X1 U4821 ( .A(n2121),  .B(n3829),  .C(n2125),  .D(n3957), .Y(n4257));
   INVX1 U4822 ( .A(w_mem_inst_w_mem[419]), .Y(n3957));
   INVX1 U4823 ( .A(w_mem_inst_w_mem[355]), .Y(n3829));
   NAND2X1 U4824 ( .A(n2119),  .B(n4085), .Y(n4256));
   INVX1 U4825 ( .A(w_mem_inst_w_mem[483]), .Y(n4085));
   NAND3X1 U4826 ( .A(n4258),  .B(n4259),  .C(n4260), .Y(n4254));
   AOI22X1 U4827 ( .A(n4158),  .B(n4021),  .C(n2123),  .D(n3701), .Y(n4260));
   INVX1 U4828 ( .A(w_mem_inst_w_mem[291]), .Y(n3701));
   INVX1 U4829 ( .A(w_mem_inst_w_mem[451]), .Y(n4021));
   NAND2X1 U4830 ( .A(n3106),  .B(n3637), .Y(n4259));
   INVX1 U4831 ( .A(w_mem_inst_w_mem[259]), .Y(n3637));
   AOI22X1 U4832 ( .A(n4160),  .B(n3765),  .C(n4161),  .D(n3893), .Y(n4258));
   INVX1 U4833 ( .A(w_mem_inst_w_mem[387]), .Y(n3893));
   INVX1 U4834 ( .A(w_mem_inst_w_mem[323]), .Y(n3765));
   NAND3X1 U4835 ( .A(n4261),  .B(n4262),  .C(n4263), .Y(n4252));
   AND2X1 U4836 ( .A(n4264),  .B(n4265), .Y(n4263));
   AOI22X1 U4837 ( .A(n4158),  .B(n3509),  .C(n2123),  .D(n3189), .Y(n4265));
   INVX1 U4838 ( .A(w_mem_inst_w_mem[35]), .Y(n3189));
   INVX1 U4839 ( .A(w_mem_inst_w_mem[195]), .Y(n3509));
   AOI22X1 U4840 ( .A(n2121),  .B(n3317),  .C(n2125),  .D(n3445), .Y(n4264));
   INVX1 U4841 ( .A(w_mem_inst_w_mem[163]), .Y(puf_10_wire_3));
   INVX1 U4842 ( .A(w_mem_inst_w_mem[99]), .Y(n3317));
   OAI21X1 U4843 ( .A(n4160),  .B(n3381),  .C(n4266), .Y(n4262));
   AOI21X1 U4844 ( .A(w_mem_inst_w_mem[67]),  .B(n2958),  .C(n4169), .Y(n4266));
   INVX1 U4845 ( .A(w_mem_inst_w_mem[131]), .Y(n3381));
   AOI22X1 U4846 ( .A(n2119),  .B(n3573),  .C(n2117),  .D(n4267), .Y(n4261));
   NAND2X1 U4847 ( .A(n4442),  .B(w_mem_inst_w_mem[3]), .Y(n4267));
   INVX1 U4848 ( .A(w_mem_inst_w_mem[227]), .Y(n3573));
   NAND3X1 U4849 ( .A(n4149),  .B(n4272),  .C(n4273), .Y(n4271));
   AOI22X1 U4850 ( .A(n2121),  .B(n3885),  .C(n2125),  .D(n4013), .Y(n4273));
   INVX1 U4851 ( .A(w_mem_inst_w_mem[447]), .Y(n4013));
   INVX1 U4852 ( .A(w_mem_inst_w_mem[383]), .Y(n3885));
   NAND2X1 U4853 ( .A(n2119),  .B(n4141), .Y(n4272));
   INVX1 U4854 ( .A(w_mem_inst_w_mem[511]), .Y(n4141));
   NAND3X1 U4855 ( .A(n4274),  .B(n4275),  .C(n4276), .Y(n4270));
   AOI22X1 U4856 ( .A(n4158),  .B(n4077),  .C(n2123),  .D(n3757), .Y(n4276));
   INVX1 U4857 ( .A(w_mem_inst_w_mem[319]), .Y(n3757));
   INVX1 U4858 ( .A(w_mem_inst_w_mem[479]), .Y(n4077));
   NAND2X1 U4859 ( .A(n3106),  .B(n3693), .Y(n4275));
   INVX1 U4860 ( .A(w_mem_inst_w_mem[287]), .Y(n3693));
   AOI22X1 U4861 ( .A(n4160),  .B(n3821),  .C(n4161),  .D(n3949), .Y(n4274));
   INVX1 U4862 ( .A(w_mem_inst_w_mem[415]), .Y(n3949));
   INVX1 U4863 ( .A(w_mem_inst_w_mem[351]), .Y(n3821));
   NAND3X1 U4864 ( .A(n4277),  .B(n4278),  .C(n4279), .Y(n4268));
   AND2X1 U4865 ( .A(n4280),  .B(n4281), .Y(n4279));
   AOI22X1 U4866 ( .A(n4158),  .B(n3565),  .C(n2123),  .D(n3245), .Y(n4281));
   INVX1 U4867 ( .A(w_mem_inst_w_mem[63]), .Y(n3245));
   INVX1 U4868 ( .A(w_mem_inst_w_mem[223]), .Y(n3565));
   AOI22X1 U4869 ( .A(n2121),  .B(n3373),  .C(n2125),  .D(n3501), .Y(n4280));
   INVX1 U4870 ( .A(w_mem_inst_w_mem[191]), .Y(n3501));
   INVX1 U4871 ( .A(w_mem_inst_w_mem[127]), .Y(n3373));
   OAI21X1 U4872 ( .A(n4160),  .B(n3437),  .C(n4282), .Y(n4278));
   AOI21X1 U4873 ( .A(w_mem_inst_w_mem[95]),  .B(n2958),  .C(n4169), .Y(n4282));
   INVX1 U4874 ( .A(w_mem_inst_w_mem[159]), .Y(n3437));
   AOI22X1 U4875 ( .A(n2119),  .B(n3629),  .C(n2117),  .D(n4283), .Y(n4277));
   NAND2X1 U4876 ( .A(n4442),  .B(w_mem_inst_w_mem[31]), .Y(n4283));
   INVX1 U4877 ( .A(w_mem_inst_w_mem[255]), .Y(n3629));
   NAND3X1 U4878 ( .A(n4149),  .B(n4288),  .C(n4289), .Y(n4287));
   AOI22X1 U4879 ( .A(n2121),  .B(n3883),  .C(n2125),  .D(n4011), .Y(n4289));
   INVX1 U4880 ( .A(w_mem_inst_w_mem[446]), .Y(n4011));
   INVX1 U4881 ( .A(w_mem_inst_w_mem[382]), .Y(n3883));
   NAND2X1 U4882 ( .A(n2119),  .B(n4139), .Y(n4288));
   INVX1 U4883 ( .A(w_mem_inst_w_mem[510]), .Y(n4139));
   NAND3X1 U4884 ( .A(n4290),  .B(n4291),  .C(n4292), .Y(n4286));
   AOI22X1 U4885 ( .A(n4158),  .B(n4075),  .C(n2123),  .D(n3755), .Y(n4292));
   INVX1 U4886 ( .A(w_mem_inst_w_mem[318]), .Y(n3755));
   INVX1 U4887 ( .A(w_mem_inst_w_mem[478]), .Y(n4075));
   NAND2X1 U4888 ( .A(n3106),  .B(n3691), .Y(n4291));
   INVX1 U4889 ( .A(w_mem_inst_w_mem[286]), .Y(n3691));
   AOI22X1 U4890 ( .A(n4160),  .B(n3819),  .C(n4161),  .D(n3947), .Y(n4290));
   INVX1 U4891 ( .A(w_mem_inst_w_mem[414]), .Y(n3947));
   INVX1 U4892 ( .A(w_mem_inst_w_mem[350]), .Y(n3819));
   NAND3X1 U4893 ( .A(n4293),  .B(n4294),  .C(n4295), .Y(n4284));
   AND2X1 U4894 ( .A(n4296),  .B(n4297), .Y(n4295));
   AOI22X1 U4895 ( .A(n4158),  .B(n3563),  .C(n2123),  .D(n3243), .Y(n4297));
   INVX1 U4896 ( .A(w_mem_inst_w_mem[62]), .Y(n3243));
   INVX1 U4897 ( .A(w_mem_inst_w_mem[222]), .Y(n3563));
   AOI22X1 U4898 ( .A(n2121),  .B(n3371),  .C(n2125),  .D(n3499), .Y(n4296));
   INVX1 U4899 ( .A(w_mem_inst_w_mem[190]), .Y(n3499));
   INVX1 U4900 ( .A(w_mem_inst_w_mem[126]), .Y(n3371));
   OAI21X1 U4901 ( .A(n4160),  .B(n3435),  .C(n4298), .Y(n4294));
   AOI21X1 U4902 ( .A(w_mem_inst_w_mem[94]),  .B(n2958),  .C(n4169), .Y(n4298));
   INVX1 U4903 ( .A(w_mem_inst_w_mem[158]), .Y(n3435));
   AOI22X1 U4904 ( .A(n2119),  .B(n3627),  .C(n2117),  .D(n4299), .Y(n4293));
   NAND2X1 U4905 ( .A(n4442),  .B(w_mem_inst_w_mem[30]), .Y(n4299));
   INVX1 U4906 ( .A(w_mem_inst_w_mem[254]), .Y(n3627));
   NAND3X1 U4907 ( .A(n4149),  .B(n4304),  .C(n4305), .Y(n4303));
   AOI22X1 U4908 ( .A(n2121),  .B(n3827),  .C(n2125),  .D(n3955), .Y(n4305));
   INVX1 U4909 ( .A(w_mem_inst_w_mem[418]), .Y(n3955));
   INVX1 U4910 ( .A(w_mem_inst_w_mem[354]), .Y(n3827));
   NAND2X1 U4911 ( .A(n2119),  .B(n4083), .Y(n4304));
   INVX1 U4912 ( .A(w_mem_inst_w_mem[482]), .Y(n4083));
   NAND3X1 U4913 ( .A(n4306),  .B(n4307),  .C(n4308), .Y(n4302));
   AOI22X1 U4914 ( .A(n4158),  .B(n4019),  .C(n2123),  .D(n3699), .Y(n4308));
   INVX1 U4915 ( .A(w_mem_inst_w_mem[290]), .Y(n3699));
   INVX1 U4916 ( .A(w_mem_inst_w_mem[450]), .Y(n4019));
   NAND2X1 U4917 ( .A(n3106),  .B(n3635), .Y(n4307));
   INVX1 U4918 ( .A(w_mem_inst_w_mem[258]), .Y(n3635));
   AOI22X1 U4919 ( .A(n4160),  .B(n3763),  .C(n4161),  .D(n3891), .Y(n4306));
   INVX1 U4920 ( .A(w_mem_inst_w_mem[386]), .Y(n3891));
   INVX1 U4921 ( .A(w_mem_inst_w_mem[322]), .Y(n3763));
   NAND3X1 U4922 ( .A(n4309),  .B(n4310),  .C(n4311), .Y(n4300));
   AND2X1 U4923 ( .A(n4312),  .B(n4313), .Y(n4311));
   AOI22X1 U4924 ( .A(n4158),  .B(n3507),  .C(n2123),  .D(n3187), .Y(n4313));
   INVX1 U4925 ( .A(w_mem_inst_w_mem[34]), .Y(n3187));
   INVX1 U4926 ( .A(w_mem_inst_w_mem[194]), .Y(n3507));
   AOI22X1 U4927 ( .A(n2121),  .B(n3315),  .C(n2125),  .D(n3443), .Y(n4312));
   INVX1 U4928 ( .A(w_mem_inst_w_mem[162]), .Y(n3443));
   INVX1 U4929 ( .A(w_mem_inst_w_mem[98]), .Y(n3315));
   OAI21X1 U4930 ( .A(n4160),  .B(n3379),  .C(n4314), .Y(n4310));
   AOI21X1 U4931 ( .A(w_mem_inst_w_mem[66]),  .B(n2958),  .C(n4169), .Y(n4314));
   INVX1 U4932 ( .A(w_mem_inst_w_mem[130]), .Y(n3379));
   AOI22X1 U4933 ( .A(n2119),  .B(n3571),  .C(n2117),  .D(n4315), .Y(n4309));
   NAND2X1 U4934 ( .A(n4442),  .B(w_mem_inst_w_mem[2]), .Y(n4315));
   INVX1 U4935 ( .A(w_mem_inst_w_mem[226]), .Y(n3571));
   NAND3X1 U4936 ( .A(n4149),  .B(n4320),  .C(n4321), .Y(n4319));
   AOI22X1 U4937 ( .A(n2121),  .B(n3881),  .C(n2125),  .D(n4009), .Y(n4321));
   INVX1 U4938 ( .A(w_mem_inst_w_mem[445]), .Y(n4009));
   INVX1 U4939 ( .A(w_mem_inst_w_mem[381]), .Y(n3881));
   NAND2X1 U4940 ( .A(n2119),  .B(n4137), .Y(n4320));
   INVX1 U4941 ( .A(w_mem_inst_w_mem[509]), .Y(n4137));
   NAND3X1 U4942 ( .A(n4322),  .B(n4323),  .C(n4324), .Y(n4318));
   AOI22X1 U4943 ( .A(n4158),  .B(n4073),  .C(n2123),  .D(n3753), .Y(n4324));
   INVX1 U4944 ( .A(w_mem_inst_w_mem[317]), .Y(n3753));
   INVX1 U4945 ( .A(w_mem_inst_w_mem[477]), .Y(n4073));
   NAND2X1 U4946 ( .A(n3106),  .B(n3689), .Y(n4323));
   INVX1 U4947 ( .A(w_mem_inst_w_mem[285]), .Y(n3689));
   AOI22X1 U4948 ( .A(n4160),  .B(n3817),  .C(n4161),  .D(n3945), .Y(n4322));
   INVX1 U4949 ( .A(w_mem_inst_w_mem[413]), .Y(n3945));
   INVX1 U4950 ( .A(w_mem_inst_w_mem[349]), .Y(n3817));
   NAND3X1 U4951 ( .A(n4325),  .B(n4326),  .C(n4327), .Y(n4316));
   AND2X1 U4952 ( .A(n4328),  .B(n4329), .Y(n4327));
   AOI22X1 U4953 ( .A(n4158),  .B(n3561),  .C(n2123),  .D(n3241), .Y(n4329));
   INVX1 U4954 ( .A(w_mem_inst_w_mem[61]), .Y(n3241));
   INVX1 U4955 ( .A(w_mem_inst_w_mem[221]), .Y(n3561));
   AOI22X1 U4956 ( .A(n2121),  .B(n3369),  .C(n2125),  .D(n3497), .Y(n4328));
   INVX1 U4957 ( .A(w_mem_inst_w_mem[189]), .Y(n3497));
   INVX1 U4958 ( .A(w_mem_inst_w_mem[125]), .Y(n3369));
   OAI21X1 U4959 ( .A(n4160),  .B(n3433),  .C(n4330), .Y(n4326));
   AOI21X1 U4960 ( .A(w_mem_inst_w_mem[93]),  .B(n2958),  .C(n4169), .Y(n4330));
   INVX1 U4961 ( .A(w_mem_inst_w_mem[157]), .Y(n3433));
   AOI22X1 U4962 ( .A(n2119),  .B(n3625),  .C(n2117),  .D(n4331), .Y(n4325));
   NAND2X1 U4963 ( .A(n4442),  .B(w_mem_inst_w_mem[29]), .Y(n4331));
   INVX1 U4964 ( .A(w_mem_inst_w_mem[253]), .Y(n3625));
   NAND3X1 U4965 ( .A(n4149),  .B(n4336),  .C(n4337), .Y(n4335));
   AOI22X1 U4966 ( .A(n2121),  .B(n3879),  .C(n2125),  .D(n4007), .Y(n4337));
   INVX1 U4967 ( .A(w_mem_inst_w_mem[444]), .Y(n4007));
   INVX1 U4968 ( .A(w_mem_inst_w_mem[380]), .Y(n3879));
   NAND2X1 U4969 ( .A(n2119),  .B(n4135), .Y(n4336));
   INVX1 U4970 ( .A(w_mem_inst_w_mem[508]), .Y(n4135));
   NAND3X1 U4971 ( .A(n4338),  .B(n4339),  .C(n4340), .Y(n4334));
   AOI22X1 U4972 ( .A(n4158),  .B(n4071),  .C(n2123),  .D(n3751), .Y(n4340));
   INVX1 U4973 ( .A(w_mem_inst_w_mem[316]), .Y(n3751));
   INVX1 U4974 ( .A(w_mem_inst_w_mem[476]), .Y(n4071));
   NAND2X1 U4975 ( .A(n3106),  .B(n3687), .Y(n4339));
   INVX1 U4976 ( .A(w_mem_inst_w_mem[284]), .Y(n3687));
   AOI22X1 U4977 ( .A(n4160),  .B(n3815),  .C(n4161),  .D(n3943), .Y(n4338));
   INVX1 U4978 ( .A(w_mem_inst_w_mem[412]), .Y(n3943));
   INVX1 U4979 ( .A(w_mem_inst_w_mem[348]), .Y(n3815));
   NAND3X1 U4980 ( .A(n4341),  .B(n4342),  .C(n4343), .Y(n4332));
   AND2X1 U4981 ( .A(n4344),  .B(n4345), .Y(n4343));
   AOI22X1 U4982 ( .A(n4158),  .B(n3559),  .C(n2123),  .D(n3239), .Y(n4345));
   INVX1 U4983 ( .A(w_mem_inst_w_mem[60]), .Y(n3239));
   INVX1 U4984 ( .A(w_mem_inst_w_mem[220]), .Y(n3559));
   AOI22X1 U4985 ( .A(n2121),  .B(n3367),  .C(n2125),  .D(n3495), .Y(n4344));
   INVX1 U4986 ( .A(w_mem_inst_w_mem[188]), .Y(n3495));
   INVX1 U4987 ( .A(w_mem_inst_w_mem[124]), .Y(n3367));
   OAI21X1 U4988 ( .A(n4160),  .B(n3431),  .C(n4346), .Y(n4342));
   AOI21X1 U4989 ( .A(w_mem_inst_w_mem[92]),  .B(n2958),  .C(n4169), .Y(n4346));
   INVX1 U4990 ( .A(w_mem_inst_w_mem[156]), .Y(n3431));
   AOI22X1 U4991 ( .A(n2119),  .B(n3623),  .C(n2117),  .D(n4347), .Y(n4341));
   NAND2X1 U4992 ( .A(n4442),  .B(w_mem_inst_w_mem[28]), .Y(n4347));
   INVX1 U4993 ( .A(w_mem_inst_w_mem[252]), .Y(n3623));
   NAND3X1 U4994 ( .A(n4149),  .B(n4352),  .C(n4353), .Y(n4351));
   AOI22X1 U4995 ( .A(n2121),  .B(n3877),  .C(n2125),  .D(n4005), .Y(n4353));
   INVX1 U4996 ( .A(w_mem_inst_w_mem[443]), .Y(n4005));
   INVX1 U4997 ( .A(w_mem_inst_w_mem[379]), .Y(n3877));
   NAND2X1 U4998 ( .A(n2119),  .B(n4133), .Y(n4352));
   INVX1 U4999 ( .A(w_mem_inst_w_mem[507]), .Y(n4133));
   NAND3X1 U5000 ( .A(n4354),  .B(n4355),  .C(n4356), .Y(n4350));
   AOI22X1 U5001 ( .A(n4158),  .B(n4069),  .C(n2123),  .D(n3749), .Y(n4356));
   INVX1 U5002 ( .A(w_mem_inst_w_mem[315]), .Y(n3749));
   INVX1 U5003 ( .A(w_mem_inst_w_mem[475]), .Y(n4069));
   NAND2X1 U5004 ( .A(n3106),  .B(n3685), .Y(n4355));
   INVX1 U5005 ( .A(w_mem_inst_w_mem[283]), .Y(n3685));
   AOI22X1 U5006 ( .A(n4160),  .B(n3813),  .C(n4161),  .D(n3941), .Y(n4354));
   INVX1 U5007 ( .A(w_mem_inst_w_mem[411]), .Y(n3941));
   INVX1 U5008 ( .A(w_mem_inst_w_mem[347]), .Y(n3813));
   NAND3X1 U5009 ( .A(n4357),  .B(n4358),  .C(n4359), .Y(n4348));
   AND2X1 U5010 ( .A(n4360),  .B(n4361), .Y(n4359));
   AOI22X1 U5011 ( .A(n4158),  .B(n3557),  .C(n2123),  .D(n3237), .Y(n4361));
   INVX1 U5012 ( .A(w_mem_inst_w_mem[59]), .Y(n3237));
   INVX1 U5013 ( .A(w_mem_inst_w_mem[219]), .Y(n3557));
   AOI22X1 U5014 ( .A(n2121),  .B(n3365),  .C(n2125),  .D(n3493), .Y(n4360));
   INVX1 U5015 ( .A(w_mem_inst_w_mem[187]), .Y(n3493));
   INVX1 U5016 ( .A(w_mem_inst_w_mem[123]), .Y(n3365));
   OAI21X1 U5017 ( .A(n4160),  .B(n3429),  .C(n4362), .Y(n4358));
   AOI21X1 U5018 ( .A(w_mem_inst_w_mem[91]),  .B(n2958),  .C(n4169), .Y(n4362));
   INVX1 U5019 ( .A(w_mem_inst_w_mem[155]), .Y(n3429));
   AOI22X1 U5020 ( .A(n2119),  .B(n3621),  .C(n2117),  .D(n4363), .Y(n4357));
   NAND2X1 U5021 ( .A(n4442),  .B(w_mem_inst_w_mem[27]), .Y(n4363));
   INVX1 U5022 ( .A(w_mem_inst_w_mem[251]), .Y(n3621));
   NAND3X1 U5023 ( .A(n4149),  .B(n4368),  .C(n4369), .Y(n4367));
   AOI22X1 U5024 ( .A(n2121),  .B(n3875),  .C(n2125),  .D(n4003), .Y(n4369));
   INVX1 U5025 ( .A(w_mem_inst_w_mem[442]), .Y(n4003));
   INVX1 U5026 ( .A(w_mem_inst_w_mem[378]), .Y(n3875));
   NAND2X1 U5027 ( .A(n2119),  .B(n4131), .Y(n4368));
   INVX1 U5028 ( .A(w_mem_inst_w_mem[506]), .Y(n4131));
   NAND3X1 U5029 ( .A(n4370),  .B(n4371),  .C(n4372), .Y(n4366));
   AOI22X1 U5030 ( .A(n4158),  .B(n4067),  .C(n2123),  .D(n3747), .Y(n4372));
   INVX1 U5031 ( .A(w_mem_inst_w_mem[314]), .Y(n3747));
   INVX1 U5032 ( .A(w_mem_inst_w_mem[474]), .Y(n4067));
   NAND2X1 U5033 ( .A(n3106),  .B(n3683), .Y(n4371));
   INVX1 U5034 ( .A(w_mem_inst_w_mem[282]), .Y(n3683));
   AOI22X1 U5035 ( .A(n4160),  .B(n3811),  .C(n4161),  .D(n3939), .Y(n4370));
   INVX1 U5036 ( .A(w_mem_inst_w_mem[410]), .Y(n3939));
   INVX1 U5037 ( .A(w_mem_inst_w_mem[346]), .Y(n3811));
   NAND3X1 U5038 ( .A(n4373),  .B(n4374),  .C(n4375), .Y(n4364));
   AND2X1 U5039 ( .A(n4376),  .B(n4377), .Y(n4375));
   AOI22X1 U5040 ( .A(n4158),  .B(n3555),  .C(n2123),  .D(n3235), .Y(n4377));
   INVX1 U5041 ( .A(w_mem_inst_w_mem[58]), .Y(n3235));
   INVX1 U5042 ( .A(w_mem_inst_w_mem[218]), .Y(n3555));
   AOI22X1 U5043 ( .A(n2121),  .B(n3363),  .C(n2125),  .D(n3491), .Y(n4376));
   INVX1 U5044 ( .A(w_mem_inst_w_mem[186]), .Y(n3491));
   INVX1 U5045 ( .A(w_mem_inst_w_mem[122]), .Y(n3363));
   OAI21X1 U5046 ( .A(n4160),  .B(n3427),  .C(n4378), .Y(n4374));
   AOI21X1 U5047 ( .A(w_mem_inst_w_mem[90]),  .B(n2958),  .C(n4169), .Y(n4378));
   INVX1 U5048 ( .A(w_mem_inst_w_mem[154]), .Y(n3427));
   AOI22X1 U5049 ( .A(n2119),  .B(n3619),  .C(n2117),  .D(n4379), .Y(n4373));
   NAND2X1 U5050 ( .A(n4442),  .B(w_mem_inst_w_mem[26]), .Y(n4379));
   INVX1 U5051 ( .A(w_mem_inst_w_mem[250]), .Y(n3619));
   NAND3X1 U5052 ( .A(n4149),  .B(n4384),  .C(n4385), .Y(n4383));
   AOI22X1 U5053 ( .A(n2121),  .B(n3873),  .C(n2125),  .D(n4001), .Y(n4385));
   INVX1 U5054 ( .A(w_mem_inst_w_mem[441]), .Y(n4001));
   INVX1 U5055 ( .A(w_mem_inst_w_mem[377]), .Y(n3873));
   NAND2X1 U5056 ( .A(n2119),  .B(n4129), .Y(n4384));
   INVX1 U5057 ( .A(w_mem_inst_w_mem[505]), .Y(n4129));
   NAND3X1 U5058 ( .A(n4386),  .B(n4387),  .C(n4388), .Y(n4382));
   AOI22X1 U5059 ( .A(n4158),  .B(n4065),  .C(n2123),  .D(n3745), .Y(n4388));
   INVX1 U5060 ( .A(w_mem_inst_w_mem[313]), .Y(n3745));
   INVX1 U5061 ( .A(w_mem_inst_w_mem[473]), .Y(n4065));
   NAND2X1 U5062 ( .A(n3106),  .B(n3681), .Y(n4387));
   INVX1 U5063 ( .A(w_mem_inst_w_mem[281]), .Y(n3681));
   AOI22X1 U5064 ( .A(n4160),  .B(n3809),  .C(n4161),  .D(n3937), .Y(n4386));
   INVX1 U5065 ( .A(w_mem_inst_w_mem[409]), .Y(n3937));
   INVX1 U5066 ( .A(w_mem_inst_w_mem[345]), .Y(n3809));
   NAND3X1 U5067 ( .A(n4389),  .B(n4390),  .C(n4391), .Y(n4380));
   AND2X1 U5068 ( .A(n4392),  .B(n4393), .Y(n4391));
   AOI22X1 U5069 ( .A(n4158),  .B(n3553),  .C(n2123),  .D(n3233), .Y(n4393));
   INVX1 U5070 ( .A(w_mem_inst_w_mem[57]), .Y(n3233));
   INVX1 U5071 ( .A(w_mem_inst_w_mem[217]), .Y(n3553));
   AOI22X1 U5072 ( .A(n2121),  .B(n3361),  .C(n2125),  .D(n3489), .Y(n4392));
   INVX1 U5073 ( .A(w_mem_inst_w_mem[185]), .Y(n3489));
   INVX1 U5074 ( .A(w_mem_inst_w_mem[121]), .Y(n3361));
   OAI21X1 U5075 ( .A(n4160),  .B(n3425),  .C(n4394), .Y(n4390));
   AOI21X1 U5076 ( .A(w_mem_inst_w_mem[89]),  .B(n2958),  .C(n4169), .Y(n4394));
   INVX1 U5077 ( .A(w_mem_inst_w_mem[153]), .Y(n3425));
   AOI22X1 U5078 ( .A(n2119),  .B(n3617),  .C(n2117),  .D(n4395), .Y(n4389));
   NAND2X1 U5079 ( .A(n4442),  .B(w_mem_inst_w_mem[25]), .Y(n4395));
   INVX1 U5080 ( .A(w_mem_inst_w_mem[249]), .Y(n3617));
   NAND3X1 U5081 ( .A(n4149),  .B(n4400),  .C(n4401), .Y(n4399));
   AOI22X1 U5082 ( .A(n2121),  .B(n3871),  .C(n2125),  .D(n3999), .Y(n4401));
   INVX1 U5083 ( .A(w_mem_inst_w_mem[440]), .Y(n3999));
   INVX1 U5084 ( .A(w_mem_inst_w_mem[376]), .Y(n3871));
   NAND2X1 U5085 ( .A(n2119),  .B(n4127), .Y(n4400));
   INVX1 U5086 ( .A(w_mem_inst_w_mem[504]), .Y(n4127));
   NAND3X1 U5087 ( .A(n4402),  .B(n4403),  .C(n4404), .Y(n4398));
   AOI22X1 U5088 ( .A(n4158),  .B(n4063),  .C(n2123),  .D(n3743), .Y(n4404));
   INVX1 U5089 ( .A(w_mem_inst_w_mem[312]), .Y(n3743));
   INVX1 U5090 ( .A(w_mem_inst_w_mem[472]), .Y(n4063));
   NAND2X1 U5091 ( .A(n3106),  .B(n3679), .Y(n4403));
   INVX1 U5092 ( .A(w_mem_inst_w_mem[280]), .Y(n3679));
   AOI22X1 U5093 ( .A(n4160),  .B(n3807),  .C(n4161),  .D(n3935), .Y(n4402));
   INVX1 U5094 ( .A(w_mem_inst_w_mem[408]), .Y(n3935));
   INVX1 U5095 ( .A(w_mem_inst_w_mem[344]), .Y(n3807));
   NAND3X1 U5096 ( .A(n4405),  .B(n4406),  .C(n4407), .Y(n4396));
   AND2X1 U5097 ( .A(n4408),  .B(n4409), .Y(n4407));
   AOI22X1 U5098 ( .A(n4158),  .B(n3551),  .C(n2123),  .D(n3231), .Y(n4409));
   INVX1 U5099 ( .A(w_mem_inst_w_mem[56]), .Y(n3231));
   INVX1 U5100 ( .A(w_mem_inst_w_mem[216]), .Y(n3551));
   AOI22X1 U5101 ( .A(n2121),  .B(n3359),  .C(n2125),  .D(n3487), .Y(n4408));
   INVX1 U5102 ( .A(w_mem_inst_w_mem[184]), .Y(n3487));
   INVX1 U5103 ( .A(w_mem_inst_w_mem[120]), .Y(n3359));
   OAI21X1 U5104 ( .A(n4160),  .B(n3423),  .C(n4410), .Y(n4406));
   AOI21X1 U5105 ( .A(w_mem_inst_w_mem[88]),  .B(n2958),  .C(n4169), .Y(n4410));
   INVX1 U5106 ( .A(w_mem_inst_w_mem[152]), .Y(n3423));
   AOI22X1 U5107 ( .A(n2119),  .B(n3615),  .C(n2117),  .D(n4411), .Y(n4405));
   NAND2X1 U5108 ( .A(n4442),  .B(w_mem_inst_w_mem[24]), .Y(n4411));
   INVX1 U5109 ( .A(w_mem_inst_w_mem[248]), .Y(n3615));
   NAND3X1 U5110 ( .A(n4149),  .B(n4416),  .C(n4417), .Y(n4415));
   AOI22X1 U5111 ( .A(n2121),  .B(n3869),  .C(n2125),  .D(n3997), .Y(n4417));
   INVX1 U5112 ( .A(w_mem_inst_w_mem[439]), .Y(n3997));
   INVX1 U5113 ( .A(w_mem_inst_w_mem[375]), .Y(n3869));
   NAND2X1 U5114 ( .A(n2119),  .B(n4125), .Y(n4416));
   INVX1 U5115 ( .A(w_mem_inst_w_mem[503]), .Y(n4125));
   NAND3X1 U5116 ( .A(n4418),  .B(n4419),  .C(n4420), .Y(n4414));
   AOI22X1 U5117 ( .A(n4158),  .B(n4061),  .C(n2123),  .D(n3741), .Y(n4420));
   INVX1 U5118 ( .A(w_mem_inst_w_mem[311]), .Y(n3741));
   INVX1 U5119 ( .A(w_mem_inst_w_mem[471]), .Y(n4061));
   NAND2X1 U5120 ( .A(n3106),  .B(n3677), .Y(n4419));
   INVX1 U5121 ( .A(w_mem_inst_w_mem[279]), .Y(n3677));
   AOI22X1 U5122 ( .A(n4160),  .B(n3805),  .C(n4161),  .D(n3933), .Y(n4418));
   INVX1 U5123 ( .A(w_mem_inst_w_mem[407]), .Y(n3933));
   INVX1 U5124 ( .A(w_mem_inst_w_mem[343]), .Y(n3805));
   NAND3X1 U5125 ( .A(n4421),  .B(n4422),  .C(n4423), .Y(n4412));
   AND2X1 U5126 ( .A(n4424),  .B(n4425), .Y(n4423));
   AOI22X1 U5127 ( .A(n4158),  .B(n3549),  .C(n2123),  .D(n3229), .Y(n4425));
   INVX1 U5128 ( .A(w_mem_inst_w_mem[55]), .Y(n3229));
   INVX1 U5129 ( .A(w_mem_inst_w_mem[215]), .Y(n3549));
   AOI22X1 U5130 ( .A(n2121),  .B(n3357),  .C(n2125),  .D(n3485), .Y(n4424));
   INVX1 U5131 ( .A(w_mem_inst_w_mem[183]), .Y(n3485));
   INVX1 U5132 ( .A(w_mem_inst_w_mem[119]), .Y(n3357));
   OAI21X1 U5133 ( .A(n4160),  .B(n3421),  .C(n4426), .Y(n4422));
   AOI21X1 U5134 ( .A(w_mem_inst_w_mem[87]),  .B(n2958),  .C(n4169), .Y(n4426));
   INVX1 U5135 ( .A(w_mem_inst_w_mem[151]), .Y(n3421));
   AOI22X1 U5136 ( .A(n2119),  .B(n3613),  .C(n2117),  .D(n4427), .Y(n4421));
   NAND2X1 U5137 ( .A(n4442),  .B(w_mem_inst_w_mem[23]), .Y(n4427));
   INVX1 U5138 ( .A(w_mem_inst_w_mem[247]), .Y(n3613));
   NAND3X1 U5139 ( .A(n4149),  .B(n4432),  .C(n4433), .Y(n4431));
   AOI22X1 U5140 ( .A(n2121),  .B(n3867),  .C(n2125),  .D(n3995), .Y(n4433));
   INVX1 U5141 ( .A(w_mem_inst_w_mem[438]), .Y(n3995));
   INVX1 U5142 ( .A(w_mem_inst_w_mem[374]), .Y(n3867));
   NAND2X1 U5143 ( .A(n2119),  .B(n4123), .Y(n4432));
   INVX1 U5144 ( .A(w_mem_inst_w_mem[502]), .Y(n4123));
   NAND3X1 U5145 ( .A(n4434),  .B(n4435),  .C(n4436), .Y(n4430));
   AOI22X1 U5146 ( .A(n4158),  .B(n4059),  .C(n2123),  .D(n3739), .Y(n4436));
   INVX1 U5147 ( .A(w_mem_inst_w_mem[310]), .Y(n3739));
   INVX1 U5148 ( .A(w_mem_inst_w_mem[470]), .Y(n4059));
   NAND2X1 U5149 ( .A(n3106),  .B(n3675), .Y(n4435));
   INVX1 U5150 ( .A(w_mem_inst_w_mem[278]), .Y(n3675));
   AOI22X1 U5151 ( .A(n4160),  .B(n3803),  .C(n4161),  .D(n3931), .Y(n4434));
   INVX1 U5152 ( .A(w_mem_inst_w_mem[406]), .Y(n3931));
   INVX1 U5153 ( .A(w_mem_inst_w_mem[342]), .Y(n3803));
   NAND3X1 U5154 ( .A(n4437),  .B(n4438),  .C(n4439), .Y(n4428));
   AND2X1 U5155 ( .A(n4440),  .B(n4441), .Y(n4439));
   AOI22X1 U5156 ( .A(n4158),  .B(n3547),  .C(n2123),  .D(n3227), .Y(n4441));
   INVX1 U5157 ( .A(w_mem_inst_w_mem[54]), .Y(n3227));
   INVX1 U5158 ( .A(w_mem_inst_w_mem[214]), .Y(n3547));
   AOI22X1 U5159 ( .A(n2121),  .B(n3355),  .C(n2125),  .D(n3483), .Y(n4440));
   INVX1 U5160 ( .A(w_mem_inst_w_mem[182]), .Y(n3483));
   INVX1 U5161 ( .A(w_mem_inst_w_mem[118]), .Y(n3355));
   OAI21X1 U5162 ( .A(n3163),  .B(n2895),  .C(n2117), .Y(n4438));
   INVX1 U5163 ( .A(w_mem_inst_w_mem[22]), .Y(n3163));
   AOI22X1 U5164 ( .A(n2119),  .B(n3611),  .C(n4443),  .D(n4444), .Y(n4437));
   NAND2X1 U5165 ( .A(w_mem_inst_w_mem[150]),  .B(n2894), .Y(n4444));
   AOI21X1 U5166 ( .A(w_mem_inst_w_mem[86]),  .B(n2958),  .C(n4169), .Y(n4443));
   INVX1 U5167 ( .A(w_mem_inst_w_mem[246]), .Y(n3611));
   NAND3X1 U5168 ( .A(n4149),  .B(n4450),  .C(n4451), .Y(n4449));
   AOI22X1 U5169 ( .A(n2121),  .B(n3865),  .C(n2125),  .D(n3993), .Y(n4451));
   INVX1 U5170 ( .A(w_mem_inst_w_mem[437]), .Y(n3993));
   INVX1 U5171 ( .A(w_mem_inst_w_mem[373]), .Y(n3865));
   NAND2X1 U5172 ( .A(n2119),  .B(n4121), .Y(n4450));
   INVX1 U5173 ( .A(w_mem_inst_w_mem[501]), .Y(n4121));
   NAND3X1 U5174 ( .A(n4452),  .B(n4453),  .C(n4454), .Y(n4448));
   AOI22X1 U5175 ( .A(n4158),  .B(n4057),  .C(n2123),  .D(n3737), .Y(n4454));
   INVX1 U5176 ( .A(w_mem_inst_w_mem[309]), .Y(n3737));
   INVX1 U5177 ( .A(w_mem_inst_w_mem[469]), .Y(n4057));
   NAND2X1 U5178 ( .A(n3106),  .B(n3673), .Y(n4453));
   INVX1 U5179 ( .A(w_mem_inst_w_mem[277]), .Y(n3673));
   AOI22X1 U5180 ( .A(n4160),  .B(n3801),  .C(n4161),  .D(n3929), .Y(n4452));
   INVX1 U5181 ( .A(w_mem_inst_w_mem[405]), .Y(n3929));
   INVX1 U5182 ( .A(w_mem_inst_w_mem[341]), .Y(n3801));
   NAND3X1 U5183 ( .A(n4455),  .B(n4456),  .C(n4457), .Y(n4446));
   AND2X1 U5184 ( .A(n4458),  .B(n4459), .Y(n4457));
   AOI22X1 U5185 ( .A(n4158),  .B(n3545),  .C(n2123),  .D(n3225), .Y(n4459));
   INVX1 U5186 ( .A(w_mem_inst_w_mem[53]), .Y(n3225));
   INVX1 U5187 ( .A(w_mem_inst_w_mem[213]), .Y(n3545));
   AOI22X1 U5188 ( .A(n2121),  .B(n3353),  .C(n2125),  .D(n3481), .Y(n4458));
   INVX1 U5189 ( .A(w_mem_inst_w_mem[181]), .Y(n3481));
   INVX1 U5190 ( .A(w_mem_inst_w_mem[117]), .Y(n3353));
   OAI21X1 U5191 ( .A(n3161),  .B(n2895),  .C(n2117), .Y(n4456));
   INVX1 U5192 ( .A(w_mem_inst_w_mem[21]), .Y(n3161));
   AOI22X1 U5193 ( .A(n2119),  .B(n3609),  .C(n4460),  .D(n4461), .Y(n4455));
   NAND2X1 U5194 ( .A(w_mem_inst_w_mem[149]),  .B(n2894), .Y(n4461));
   AOI21X1 U5195 ( .A(w_mem_inst_w_mem[85]),  .B(n2958),  .C(n4169), .Y(n4460));
   INVX1 U5196 ( .A(w_mem_inst_w_mem[245]), .Y(n3609));
   NAND3X1 U5197 ( .A(n4149),  .B(n4466),  .C(n4467), .Y(n4465));
   AOI22X1 U5198 ( .A(n2121),  .B(n3863),  .C(n2125),  .D(n3991), .Y(n4467));
   INVX1 U5199 ( .A(w_mem_inst_w_mem[436]), .Y(n3991));
   INVX1 U5200 ( .A(w_mem_inst_w_mem[372]), .Y(n3863));
   NAND2X1 U5201 ( .A(n2119),  .B(n4119), .Y(n4466));
   INVX1 U5202 ( .A(w_mem_inst_w_mem[500]), .Y(n4119));
   NAND3X1 U5203 ( .A(n4468),  .B(n4469),  .C(n4470), .Y(n4464));
   AOI22X1 U5204 ( .A(n4158),  .B(n4055),  .C(n2123),  .D(n3735), .Y(n4470));
   INVX1 U5205 ( .A(w_mem_inst_w_mem[308]), .Y(n3735));
   INVX1 U5206 ( .A(w_mem_inst_w_mem[468]), .Y(n4055));
   NAND2X1 U5207 ( .A(n3106),  .B(n3671), .Y(n4469));
   INVX1 U5208 ( .A(w_mem_inst_w_mem[276]), .Y(n3671));
   AOI22X1 U5209 ( .A(n4160),  .B(n3799),  .C(n4161),  .D(n3927), .Y(n4468));
   INVX1 U5210 ( .A(w_mem_inst_w_mem[404]), .Y(n3927));
   INVX1 U5211 ( .A(w_mem_inst_w_mem[340]), .Y(n3799));
   NAND3X1 U5212 ( .A(n4471),  .B(n4472),  .C(n4473), .Y(n4462));
   AND2X1 U5213 ( .A(n4474),  .B(n4475), .Y(n4473));
   AOI22X1 U5214 ( .A(n4158),  .B(n3543),  .C(n2123),  .D(n3223), .Y(n4475));
   INVX1 U5215 ( .A(w_mem_inst_w_mem[52]), .Y(n3223));
   INVX1 U5216 ( .A(w_mem_inst_w_mem[212]), .Y(n3543));
   AOI22X1 U5217 ( .A(n2121),  .B(n3351),  .C(n2125),  .D(n3479), .Y(n4474));
   INVX1 U5218 ( .A(w_mem_inst_w_mem[180]), .Y(n3479));
   INVX1 U5219 ( .A(w_mem_inst_w_mem[116]), .Y(n3351));
   OAI21X1 U5220 ( .A(n3159),  .B(n2895),  .C(n2117), .Y(n4472));
   INVX1 U5221 ( .A(w_mem_inst_w_mem[20]), .Y(n3159));
   AOI22X1 U5222 ( .A(n2119),  .B(n3607),  .C(n4476),  .D(n4477), .Y(n4471));
   NAND2X1 U5223 ( .A(w_mem_inst_w_mem[148]),  .B(n2894), .Y(n4477));
   AOI21X1 U5224 ( .A(w_mem_inst_w_mem[84]),  .B(n2958),  .C(n4169), .Y(n4476));
   INVX1 U5225 ( .A(w_mem_inst_w_mem[244]), .Y(n3607));
   NAND3X1 U5226 ( .A(n4149),  .B(n4482),  .C(n4483), .Y(n4481));
   AOI22X1 U5227 ( .A(n2121),  .B(n3825),  .C(n2125),  .D(n3953), .Y(n4483));
   INVX1 U5228 ( .A(w_mem_inst_w_mem[417]), .Y(n3953));
   INVX1 U5229 ( .A(w_mem_inst_w_mem[353]), .Y(n3825));
   NAND2X1 U5230 ( .A(n2119),  .B(n4081), .Y(n4482));
   INVX1 U5231 ( .A(w_mem_inst_w_mem[481]), .Y(n4081));
   NAND3X1 U5232 ( .A(n4484),  .B(n4485),  .C(n4486), .Y(n4480));
   AOI22X1 U5233 ( .A(n4158),  .B(n4017),  .C(n2123),  .D(n3697), .Y(n4486));
   INVX1 U5234 ( .A(w_mem_inst_w_mem[289]), .Y(n3697));
   INVX1 U5235 ( .A(w_mem_inst_w_mem[449]), .Y(n4017));
   NAND2X1 U5236 ( .A(n3106),  .B(n3633), .Y(n4485));
   INVX1 U5237 ( .A(w_mem_inst_w_mem[257]), .Y(n3633));
   AOI22X1 U5238 ( .A(n4160),  .B(n3761),  .C(n4161),  .D(n3889), .Y(n4484));
   INVX1 U5239 ( .A(w_mem_inst_w_mem[385]), .Y(n3889));
   INVX1 U5240 ( .A(w_mem_inst_w_mem[321]), .Y(n3761));
   NAND3X1 U5241 ( .A(n4487),  .B(n4488),  .C(n4489), .Y(n4478));
   AND2X1 U5242 ( .A(n4490),  .B(n4491), .Y(n4489));
   AOI22X1 U5243 ( .A(n4158),  .B(n3505),  .C(n2123),  .D(n3185), .Y(n4491));
   INVX1 U5244 ( .A(w_mem_inst_w_mem[33]), .Y(n3185));
   INVX1 U5245 ( .A(w_mem_inst_w_mem[193]), .Y(n3505));
   AOI22X1 U5246 ( .A(n2121),  .B(n3313),  .C(n2125),  .D(n3441), .Y(n4490));
   INVX1 U5247 ( .A(w_mem_inst_w_mem[161]), .Y(n3441));
   INVX1 U5248 ( .A(w_mem_inst_w_mem[97]), .Y(n3313));
   OAI21X1 U5249 ( .A(n3121),  .B(n2895),  .C(n2117), .Y(n4488));
   INVX1 U5250 ( .A(w_mem_inst_w_mem[1]), .Y(n3121));
   AOI22X1 U5251 ( .A(n2119),  .B(n3569),  .C(n4492),  .D(n4493), .Y(n4487));
   NAND2X1 U5252 ( .A(w_mem_inst_w_mem[129]),  .B(n2894), .Y(n4493));
   AOI21X1 U5253 ( .A(w_mem_inst_w_mem[65]),  .B(n2958),  .C(n4169), .Y(n4492));
   INVX1 U5254 ( .A(w_mem_inst_w_mem[225]), .Y(n3569));
   NAND3X1 U5255 ( .A(n4149),  .B(n4498),  .C(n4499), .Y(n4497));
   AOI22X1 U5256 ( .A(n2121),  .B(n3861),  .C(n2125),  .D(n3989), .Y(n4499));
   INVX1 U5257 ( .A(w_mem_inst_w_mem[435]), .Y(n3989));
   INVX1 U5258 ( .A(w_mem_inst_w_mem[371]), .Y(n3861));
   NAND2X1 U5259 ( .A(n2119),  .B(n4117), .Y(n4498));
   INVX1 U5260 ( .A(w_mem_inst_w_mem[499]), .Y(n4117));
   NAND3X1 U5261 ( .A(n4500),  .B(n4501),  .C(n4502), .Y(n4496));
   AOI22X1 U5262 ( .A(n4158),  .B(n4053),  .C(n2123),  .D(n3733), .Y(n4502));
   INVX1 U5263 ( .A(w_mem_inst_w_mem[307]), .Y(n3733));
   INVX1 U5264 ( .A(w_mem_inst_w_mem[467]), .Y(n4053));
   NAND2X1 U5265 ( .A(n3106),  .B(n3669), .Y(n4501));
   INVX1 U5266 ( .A(w_mem_inst_w_mem[275]), .Y(n3669));
   AOI22X1 U5267 ( .A(n4160),  .B(n3797),  .C(n4161),  .D(n3925), .Y(n4500));
   INVX1 U5268 ( .A(w_mem_inst_w_mem[403]), .Y(n3925));
   INVX1 U5269 ( .A(w_mem_inst_w_mem[339]), .Y(n3797));
   NAND3X1 U5270 ( .A(n4503),  .B(n4504),  .C(n4505), .Y(n4494));
   AND2X1 U5271 ( .A(n4506),  .B(n4507), .Y(n4505));
   AOI22X1 U5272 ( .A(n4158),  .B(n3541),  .C(n2123),  .D(n3221), .Y(n4507));
   INVX1 U5273 ( .A(w_mem_inst_w_mem[51]), .Y(n3221));
   INVX1 U5274 ( .A(w_mem_inst_w_mem[211]), .Y(n3541));
   AOI22X1 U5275 ( .A(n2121),  .B(n3349),  .C(n2125),  .D(n3477), .Y(n4506));
   INVX1 U5276 ( .A(w_mem_inst_w_mem[179]), .Y(n3477));
   INVX1 U5277 ( .A(w_mem_inst_w_mem[115]), .Y(n3349));
   OAI21X1 U5278 ( .A(n3157),  .B(n2895),  .C(n2117), .Y(n4504));
   INVX1 U5279 ( .A(w_mem_inst_w_mem[19]), .Y(n3157));
   AOI22X1 U5280 ( .A(n2119),  .B(n3605),  .C(n4508),  .D(n4509), .Y(n4503));
   NAND2X1 U5281 ( .A(w_mem_inst_w_mem[147]),  .B(n2894), .Y(n4509));
   AOI21X1 U5282 ( .A(w_mem_inst_w_mem[83]),  .B(n2958),  .C(n4169), .Y(n4508));
   INVX1 U5283 ( .A(w_mem_inst_w_mem[243]), .Y(n3605));
   NAND3X1 U5284 ( .A(n4149),  .B(n4514),  .C(n4515), .Y(n4513));
   AOI22X1 U5285 ( .A(n2121),  .B(n3859),  .C(n2125),  .D(n3987), .Y(n4515));
   INVX1 U5286 ( .A(w_mem_inst_w_mem[434]), .Y(n3987));
   INVX1 U5287 ( .A(w_mem_inst_w_mem[370]), .Y(n3859));
   NAND2X1 U5288 ( .A(n2119),  .B(n4115), .Y(n4514));
   INVX1 U5289 ( .A(w_mem_inst_w_mem[498]), .Y(n4115));
   NAND3X1 U5290 ( .A(n4516),  .B(n4517),  .C(n4518), .Y(n4512));
   AOI22X1 U5291 ( .A(n4158),  .B(n4051),  .C(n2123),  .D(n3731), .Y(n4518));
   INVX1 U5292 ( .A(w_mem_inst_w_mem[306]), .Y(n3731));
   INVX1 U5293 ( .A(w_mem_inst_w_mem[466]), .Y(n4051));
   NAND2X1 U5294 ( .A(n3106),  .B(n3667), .Y(n4517));
   INVX1 U5295 ( .A(w_mem_inst_w_mem[274]), .Y(n3667));
   AOI22X1 U5296 ( .A(n4160),  .B(n3795),  .C(n4161),  .D(n3923), .Y(n4516));
   INVX1 U5297 ( .A(w_mem_inst_w_mem[402]), .Y(n3923));
   INVX1 U5298 ( .A(w_mem_inst_w_mem[338]), .Y(n3795));
   NAND3X1 U5299 ( .A(n4519),  .B(n4520),  .C(n4521), .Y(n4510));
   AND2X1 U5300 ( .A(n4522),  .B(n4523), .Y(n4521));
   AOI22X1 U5301 ( .A(n4158),  .B(n3539),  .C(n2123),  .D(n3219), .Y(n4523));
   INVX1 U5302 ( .A(w_mem_inst_w_mem[50]), .Y(n3219));
   INVX1 U5303 ( .A(w_mem_inst_w_mem[210]), .Y(n3539));
   AOI22X1 U5304 ( .A(n2121),  .B(n3347),  .C(n2125),  .D(n3475), .Y(n4522));
   INVX1 U5305 ( .A(w_mem_inst_w_mem[178]), .Y(n3475));
   INVX1 U5306 ( .A(w_mem_inst_w_mem[114]), .Y(n3347));
   OAI21X1 U5307 ( .A(n3155),  .B(n2895),  .C(n2117), .Y(n4520));
   INVX1 U5308 ( .A(w_mem_inst_w_mem[18]), .Y(n3155));
   AOI22X1 U5309 ( .A(n2119),  .B(n3603),  .C(n4524),  .D(n4525), .Y(n4519));
   NAND2X1 U5310 ( .A(w_mem_inst_w_mem[146]),  .B(n2894), .Y(n4525));
   AOI21X1 U5311 ( .A(w_mem_inst_w_mem[82]),  .B(n2958),  .C(n4169), .Y(n4524));
   INVX1 U5312 ( .A(w_mem_inst_w_mem[242]), .Y(n3603));
   NAND3X1 U5313 ( .A(n4149),  .B(n4530),  .C(n4531), .Y(n4529));
   AOI22X1 U5314 ( .A(n2121),  .B(n3857),  .C(n2125),  .D(n3985), .Y(n4531));
   INVX1 U5315 ( .A(w_mem_inst_w_mem[433]), .Y(n3985));
   INVX1 U5316 ( .A(w_mem_inst_w_mem[369]), .Y(n3857));
   NAND2X1 U5317 ( .A(n2119),  .B(n4113), .Y(n4530));
   INVX1 U5318 ( .A(w_mem_inst_w_mem[497]), .Y(n4113));
   NAND3X1 U5319 ( .A(n4532),  .B(n4533),  .C(n4534), .Y(n4528));
   AOI22X1 U5320 ( .A(n4158),  .B(n4049),  .C(n2123),  .D(n3729), .Y(n4534));
   INVX1 U5321 ( .A(w_mem_inst_w_mem[305]), .Y(n3729));
   INVX1 U5322 ( .A(w_mem_inst_w_mem[465]), .Y(n4049));
   NAND2X1 U5323 ( .A(n3106),  .B(n3665), .Y(n4533));
   INVX1 U5324 ( .A(w_mem_inst_w_mem[273]), .Y(n3665));
   AOI22X1 U5325 ( .A(n4160),  .B(n3793),  .C(n4161),  .D(n3921), .Y(n4532));
   INVX1 U5326 ( .A(w_mem_inst_w_mem[401]), .Y(n3921));
   INVX1 U5327 ( .A(w_mem_inst_w_mem[337]), .Y(n3793));
   NAND3X1 U5328 ( .A(n4535),  .B(n4536),  .C(n4537), .Y(n4526));
   AND2X1 U5329 ( .A(n4538),  .B(n4539), .Y(n4537));
   AOI22X1 U5330 ( .A(n4158),  .B(n3537),  .C(n2123),  .D(n3217), .Y(n4539));
   INVX1 U5331 ( .A(w_mem_inst_w_mem[49]), .Y(n3217));
   INVX1 U5332 ( .A(w_mem_inst_w_mem[209]), .Y(n3537));
   AOI22X1 U5333 ( .A(n2121),  .B(n3345),  .C(n2125),  .D(n3473), .Y(n4538));
   INVX1 U5334 ( .A(w_mem_inst_w_mem[177]), .Y(n3473));
   INVX1 U5335 ( .A(w_mem_inst_w_mem[113]), .Y(n3345));
   OAI21X1 U5336 ( .A(n3153),  .B(n2895),  .C(n2117), .Y(n4536));
   INVX1 U5337 ( .A(w_mem_inst_w_mem[17]), .Y(n3153));
   AOI22X1 U5338 ( .A(n2119),  .B(n3601),  .C(n4540),  .D(n4541), .Y(n4535));
   NAND2X1 U5339 ( .A(w_mem_inst_w_mem[145]),  .B(n2894), .Y(n4541));
   AOI21X1 U5340 ( .A(w_mem_inst_w_mem[81]),  .B(n2958),  .C(n4169), .Y(n4540));
   INVX1 U5341 ( .A(w_mem_inst_w_mem[241]), .Y(n3601));
   NAND3X1 U5342 ( .A(n4149),  .B(n4546),  .C(n4547), .Y(n4545));
   AOI22X1 U5343 ( .A(n2121),  .B(n3855),  .C(n2125),  .D(n3983), .Y(n4547));
   INVX1 U5344 ( .A(w_mem_inst_w_mem[432]), .Y(n3983));
   INVX1 U5345 ( .A(w_mem_inst_w_mem[368]), .Y(n3855));
   NAND2X1 U5346 ( .A(n2119),  .B(n4111), .Y(n4546));
   INVX1 U5347 ( .A(w_mem_inst_w_mem[496]), .Y(n4111));
   NAND3X1 U5348 ( .A(n4548),  .B(n4549),  .C(n4550), .Y(n4544));
   AOI22X1 U5349 ( .A(n4158),  .B(n4047),  .C(n2123),  .D(n3727), .Y(n4550));
   INVX1 U5350 ( .A(w_mem_inst_w_mem[304]), .Y(n3727));
   INVX1 U5351 ( .A(w_mem_inst_w_mem[464]), .Y(n4047));
   NAND2X1 U5352 ( .A(n3106),  .B(n3663), .Y(n4549));
   INVX1 U5353 ( .A(w_mem_inst_w_mem[272]), .Y(n3663));
   AOI22X1 U5354 ( .A(n4160),  .B(n3791),  .C(n4161),  .D(n3919), .Y(n4548));
   INVX1 U5355 ( .A(w_mem_inst_w_mem[400]), .Y(n3919));
   INVX1 U5356 ( .A(w_mem_inst_w_mem[336]), .Y(n3791));
   NAND3X1 U5357 ( .A(n4551),  .B(n4552),  .C(n4553), .Y(n4542));
   AND2X1 U5358 ( .A(n4554),  .B(n4555), .Y(n4553));
   AOI22X1 U5359 ( .A(n4158),  .B(n3535),  .C(n2123),  .D(n3215), .Y(n4555));
   INVX1 U5360 ( .A(w_mem_inst_w_mem[48]), .Y(n3215));
   INVX1 U5361 ( .A(w_mem_inst_w_mem[208]), .Y(n3535));
   AOI22X1 U5362 ( .A(n2121),  .B(n3343),  .C(n2125),  .D(n3471), .Y(n4554));
   INVX1 U5363 ( .A(w_mem_inst_w_mem[176]), .Y(n3471));
   INVX1 U5364 ( .A(w_mem_inst_w_mem[112]), .Y(n3343));
   OAI21X1 U5365 ( .A(n3151),  .B(n2895),  .C(n2117), .Y(n4552));
   INVX1 U5366 ( .A(w_mem_inst_w_mem[16]), .Y(n3151));
   AOI22X1 U5367 ( .A(n2119),  .B(n3599),  .C(n4556),  .D(n4557), .Y(n4551));
   NAND2X1 U5368 ( .A(w_mem_inst_w_mem[144]),  .B(n2894), .Y(n4557));
   AOI21X1 U5369 ( .A(w_mem_inst_w_mem[80]),  .B(n2958),  .C(n4169), .Y(n4556));
   INVX1 U5370 ( .A(w_mem_inst_w_mem[240]), .Y(n3599));
   NAND3X1 U5371 ( .A(n4149),  .B(n4562),  .C(n4563), .Y(n4561));
   AOI22X1 U5372 ( .A(n2121),  .B(n3853),  .C(n2125),  .D(n3981), .Y(n4563));
   INVX1 U5373 ( .A(w_mem_inst_w_mem[431]), .Y(n3981));
   INVX1 U5374 ( .A(w_mem_inst_w_mem[367]), .Y(n3853));
   NAND2X1 U5375 ( .A(n2119),  .B(n4109), .Y(n4562));
   INVX1 U5376 ( .A(w_mem_inst_w_mem[495]), .Y(n4109));
   NAND3X1 U5377 ( .A(n4564),  .B(n4565),  .C(n4566), .Y(n4560));
   AOI22X1 U5378 ( .A(n4158),  .B(n4045),  .C(n2123),  .D(n3725), .Y(n4566));
   INVX1 U5379 ( .A(w_mem_inst_w_mem[303]), .Y(n3725));
   INVX1 U5380 ( .A(w_mem_inst_w_mem[463]), .Y(n4045));
   NAND2X1 U5381 ( .A(n3106),  .B(n3661), .Y(n4565));
   INVX1 U5382 ( .A(w_mem_inst_w_mem[271]), .Y(n3661));
   AOI22X1 U5383 ( .A(n4160),  .B(n3789),  .C(n4161),  .D(n3917), .Y(n4564));
   INVX1 U5384 ( .A(w_mem_inst_w_mem[399]), .Y(n3917));
   INVX1 U5385 ( .A(w_mem_inst_w_mem[335]), .Y(n3789));
   NAND3X1 U5386 ( .A(n4567),  .B(n4568),  .C(n4569), .Y(n4558));
   AND2X1 U5387 ( .A(n4570),  .B(n4571), .Y(n4569));
   AOI22X1 U5388 ( .A(n4158),  .B(n3533),  .C(n2123),  .D(n3213), .Y(n4571));
   INVX1 U5389 ( .A(w_mem_inst_w_mem[47]), .Y(n3213));
   INVX1 U5390 ( .A(w_mem_inst_w_mem[207]), .Y(n3533));
   AOI22X1 U5391 ( .A(n2121),  .B(n3341),  .C(n2125),  .D(n3469), .Y(n4570));
   INVX1 U5392 ( .A(w_mem_inst_w_mem[175]), .Y(n3469));
   INVX1 U5393 ( .A(w_mem_inst_w_mem[111]), .Y(n3341));
   OAI21X1 U5394 ( .A(n3149),  .B(n2895),  .C(n2117), .Y(n4568));
   INVX1 U5395 ( .A(w_mem_inst_w_mem[15]), .Y(n3149));
   AOI22X1 U5396 ( .A(n2119),  .B(n3597),  .C(n4572),  .D(n4573), .Y(n4567));
   NAND2X1 U5397 ( .A(w_mem_inst_w_mem[143]),  .B(n2894), .Y(n4573));
   AOI21X1 U5398 ( .A(w_mem_inst_w_mem[79]),  .B(n2958),  .C(n4169), .Y(n4572));
   INVX1 U5399 ( .A(w_mem_inst_w_mem[239]), .Y(n3597));
   NAND3X1 U5400 ( .A(n4149),  .B(n4578),  .C(n4579), .Y(n4577));
   AOI22X1 U5401 ( .A(n2121),  .B(n3851),  .C(n2125),  .D(n3979), .Y(n4579));
   INVX1 U5402 ( .A(w_mem_inst_w_mem[430]), .Y(n3979));
   INVX1 U5403 ( .A(w_mem_inst_w_mem[366]), .Y(n3851));
   NAND2X1 U5404 ( .A(n2119),  .B(n4107), .Y(n4578));
   INVX1 U5405 ( .A(w_mem_inst_w_mem[494]), .Y(n4107));
   NAND3X1 U5406 ( .A(n4580),  .B(n4581),  .C(n4582), .Y(n4576));
   AOI22X1 U5407 ( .A(n4158),  .B(n4043),  .C(n2123),  .D(n3723), .Y(n4582));
   INVX1 U5408 ( .A(w_mem_inst_w_mem[302]), .Y(n3723));
   INVX1 U5409 ( .A(w_mem_inst_w_mem[462]), .Y(n4043));
   NAND2X1 U5410 ( .A(n3106),  .B(n3659), .Y(n4581));
   INVX1 U5411 ( .A(w_mem_inst_w_mem[270]), .Y(n3659));
   AOI22X1 U5412 ( .A(n4160),  .B(n3787),  .C(n4161),  .D(n3915), .Y(n4580));
   INVX1 U5413 ( .A(w_mem_inst_w_mem[398]), .Y(n3915));
   INVX1 U5414 ( .A(w_mem_inst_w_mem[334]), .Y(n3787));
   NAND3X1 U5415 ( .A(n4583),  .B(n4584),  .C(n4585), .Y(n4574));
   AND2X1 U5416 ( .A(n4586),  .B(n4587), .Y(n4585));
   AOI22X1 U5417 ( .A(n4158),  .B(n3531),  .C(n2123),  .D(n3211), .Y(n4587));
   INVX1 U5418 ( .A(w_mem_inst_w_mem[46]), .Y(n3211));
   INVX1 U5419 ( .A(w_mem_inst_w_mem[206]), .Y(n3531));
   AOI22X1 U5420 ( .A(n2121),  .B(n3339),  .C(n2125),  .D(n3467), .Y(n4586));
   INVX1 U5421 ( .A(w_mem_inst_w_mem[174]), .Y(n3467));
   INVX1 U5422 ( .A(w_mem_inst_w_mem[110]), .Y(n3339));
   OAI21X1 U5423 ( .A(n3147),  .B(n2895),  .C(n2117), .Y(n4584));
   INVX1 U5424 ( .A(w_mem_inst_w_mem[14]), .Y(n3147));
   AOI22X1 U5425 ( .A(n2119),  .B(n3595),  .C(n4588),  .D(n4589), .Y(n4583));
   NAND2X1 U5426 ( .A(w_mem_inst_w_mem[142]),  .B(n2894), .Y(n4589));
   AOI21X1 U5427 ( .A(w_mem_inst_w_mem[78]),  .B(n2958),  .C(n4169), .Y(n4588));
   INVX1 U5428 ( .A(w_mem_inst_w_mem[238]), .Y(n3595));
   NAND3X1 U5429 ( .A(n4149),  .B(n4594),  .C(n4595), .Y(n4593));
   AOI22X1 U5430 ( .A(n2121),  .B(n3849),  .C(n2125),  .D(n3977), .Y(n4595));
   INVX1 U5431 ( .A(w_mem_inst_w_mem[429]), .Y(n3977));
   INVX1 U5432 ( .A(w_mem_inst_w_mem[365]), .Y(n3849));
   NAND2X1 U5433 ( .A(n2119),  .B(n4105), .Y(n4594));
   INVX1 U5434 ( .A(w_mem_inst_w_mem[493]), .Y(n4105));
   NAND3X1 U5435 ( .A(n4596),  .B(n4597),  .C(n4598), .Y(n4592));
   AOI22X1 U5436 ( .A(n4158),  .B(n4041),  .C(n2123),  .D(n3721), .Y(n4598));
   INVX1 U5437 ( .A(w_mem_inst_w_mem[301]), .Y(n3721));
   INVX1 U5438 ( .A(w_mem_inst_w_mem[461]), .Y(n4041));
   NAND2X1 U5439 ( .A(n3106),  .B(n3657), .Y(n4597));
   INVX1 U5440 ( .A(w_mem_inst_w_mem[269]), .Y(n3657));
   AOI22X1 U5441 ( .A(n4160),  .B(n3785),  .C(n4161),  .D(n3913), .Y(n4596));
   INVX1 U5442 ( .A(w_mem_inst_w_mem[397]), .Y(n3913));
   INVX1 U5443 ( .A(w_mem_inst_w_mem[333]), .Y(n3785));
   NAND3X1 U5444 ( .A(n4599),  .B(n4600),  .C(n4601), .Y(n4590));
   AND2X1 U5445 ( .A(n4602),  .B(n4603), .Y(n4601));
   AOI22X1 U5446 ( .A(n4158),  .B(n3529),  .C(n2123),  .D(n3209), .Y(n4603));
   INVX1 U5447 ( .A(w_mem_inst_w_mem[45]), .Y(n3209));
   INVX1 U5448 ( .A(w_mem_inst_w_mem[205]), .Y(n3529));
   AOI22X1 U5449 ( .A(n2121),  .B(n3337),  .C(n2125),  .D(n3465), .Y(n4602));
   INVX1 U5450 ( .A(w_mem_inst_w_mem[173]), .Y(n3465));
   INVX1 U5451 ( .A(w_mem_inst_w_mem[109]), .Y(n3337));
   OAI21X1 U5452 ( .A(n3145),  .B(n2895),  .C(n2117), .Y(n4600));
   INVX1 U5453 ( .A(w_mem_inst_w_mem[13]), .Y(n3145));
   AOI22X1 U5454 ( .A(n2119),  .B(n3593),  .C(n4604),  .D(n4605), .Y(n4599));
   NAND2X1 U5455 ( .A(w_mem_inst_w_mem[141]),  .B(n2894), .Y(n4605));
   AOI21X1 U5456 ( .A(w_mem_inst_w_mem[77]),  .B(n2958),  .C(n4169), .Y(n4604));
   INVX1 U5457 ( .A(w_mem_inst_w_mem[237]), .Y(n3593));
   NAND3X1 U5458 ( .A(n4149),  .B(n4610),  .C(n4611), .Y(n4609));
   AOI22X1 U5459 ( .A(n2121),  .B(n3847),  .C(n2125),  .D(n3975), .Y(n4611));
   INVX1 U5460 ( .A(w_mem_inst_w_mem[428]), .Y(n3975));
   INVX1 U5461 ( .A(w_mem_inst_w_mem[364]), .Y(n3847));
   NAND2X1 U5462 ( .A(n2119),  .B(n4103), .Y(n4610));
   INVX1 U5463 ( .A(w_mem_inst_w_mem[492]), .Y(n4103));
   NAND3X1 U5464 ( .A(n4612),  .B(n4613),  .C(n4614), .Y(n4608));
   AOI22X1 U5465 ( .A(n4158),  .B(n4039),  .C(n2123),  .D(n3719), .Y(n4614));
   INVX1 U5466 ( .A(w_mem_inst_w_mem[300]), .Y(n3719));
   INVX1 U5467 ( .A(w_mem_inst_w_mem[460]), .Y(n4039));
   NAND2X1 U5468 ( .A(n3106),  .B(n3655), .Y(n4613));
   INVX1 U5469 ( .A(w_mem_inst_w_mem[268]), .Y(n3655));
   AOI22X1 U5470 ( .A(n4160),  .B(n3783),  .C(n4161),  .D(n3911), .Y(n4612));
   INVX1 U5471 ( .A(w_mem_inst_w_mem[396]), .Y(n3911));
   INVX1 U5472 ( .A(w_mem_inst_w_mem[332]), .Y(n3783));
   NAND3X1 U5473 ( .A(n4615),  .B(n4616),  .C(n4617), .Y(n4606));
   AND2X1 U5474 ( .A(n4618),  .B(n4619), .Y(n4617));
   AOI22X1 U5475 ( .A(n4158),  .B(n3527),  .C(n2123),  .D(n3207), .Y(n4619));
   INVX1 U5476 ( .A(w_mem_inst_w_mem[44]), .Y(n3207));
   INVX1 U5477 ( .A(w_mem_inst_w_mem[204]), .Y(n3527));
   AOI22X1 U5478 ( .A(n2121),  .B(n3335),  .C(n2125),  .D(n3463), .Y(n4618));
   INVX1 U5479 ( .A(w_mem_inst_w_mem[172]), .Y(n3463));
   INVX1 U5480 ( .A(w_mem_inst_w_mem[108]), .Y(n3335));
   OAI21X1 U5481 ( .A(n3143),  .B(n2895),  .C(n2117), .Y(n4616));
   INVX1 U5482 ( .A(w_mem_inst_w_mem[12]), .Y(n3143));
   AOI22X1 U5483 ( .A(n2119),  .B(n3591),  .C(n4620),  .D(n4621), .Y(n4615));
   NAND2X1 U5484 ( .A(w_mem_inst_w_mem[140]),  .B(n2894), .Y(n4621));
   AOI21X1 U5485 ( .A(w_mem_inst_w_mem[76]),  .B(n2958),  .C(n4169), .Y(n4620));
   INVX1 U5486 ( .A(w_mem_inst_w_mem[236]), .Y(n3591));
   NAND3X1 U5487 ( .A(n4149),  .B(n4626),  .C(n4627), .Y(n4625));
   AOI22X1 U5488 ( .A(n2121),  .B(n3845),  .C(n2125),  .D(n3973), .Y(n4627));
   INVX1 U5489 ( .A(w_mem_inst_w_mem[427]), .Y(n3973));
   INVX1 U5490 ( .A(w_mem_inst_w_mem[363]), .Y(n3845));
   NAND2X1 U5491 ( .A(n2119),  .B(n4101), .Y(n4626));
   INVX1 U5492 ( .A(w_mem_inst_w_mem[491]), .Y(n4101));
   NAND3X1 U5493 ( .A(n4628),  .B(n4629),  .C(n4630), .Y(n4624));
   AOI22X1 U5494 ( .A(n4158),  .B(n4037),  .C(n2123),  .D(n3717), .Y(n4630));
   INVX1 U5495 ( .A(w_mem_inst_w_mem[299]), .Y(n3717));
   INVX1 U5496 ( .A(w_mem_inst_w_mem[459]), .Y(n4037));
   NAND2X1 U5497 ( .A(n3106),  .B(n3653), .Y(n4629));
   INVX1 U5498 ( .A(w_mem_inst_w_mem[267]), .Y(n3653));
   AOI22X1 U5499 ( .A(n4160),  .B(n3781),  .C(n4161),  .D(n3909), .Y(n4628));
   INVX1 U5500 ( .A(w_mem_inst_w_mem[395]), .Y(n3909));
   INVX1 U5501 ( .A(w_mem_inst_w_mem[331]), .Y(n3781));
   NAND3X1 U5502 ( .A(n4631),  .B(n4632),  .C(n4633), .Y(n4622));
   AND2X1 U5503 ( .A(n4634),  .B(n4635), .Y(n4633));
   AOI22X1 U5504 ( .A(n4158),  .B(n3525),  .C(n2123),  .D(n3205), .Y(n4635));
   INVX1 U5505 ( .A(w_mem_inst_w_mem[43]), .Y(n3205));
   INVX1 U5506 ( .A(w_mem_inst_w_mem[203]), .Y(n3525));
   AOI22X1 U5507 ( .A(n2121),  .B(n3333),  .C(n2125),  .D(n3461), .Y(n4634));
   INVX1 U5508 ( .A(w_mem_inst_w_mem[171]), .Y(n3461));
   INVX1 U5509 ( .A(w_mem_inst_w_mem[107]), .Y(n3333));
   OAI21X1 U5510 ( .A(n3141),  .B(n2895),  .C(n2117), .Y(n4632));
   INVX1 U5511 ( .A(w_mem_inst_w_mem[11]), .Y(n3141));
   AOI22X1 U5512 ( .A(n2119),  .B(n3589),  .C(n4636),  .D(n4637), .Y(n4631));
   NAND2X1 U5513 ( .A(w_mem_inst_w_mem[139]),  .B(n2894), .Y(n4637));
   AOI21X1 U5514 ( .A(w_mem_inst_w_mem[75]),  .B(n2958),  .C(n4169), .Y(n4636));
   INVX1 U5515 ( .A(w_mem_inst_w_mem[235]), .Y(n3589));
   NAND3X1 U5516 ( .A(n4149),  .B(n4642),  .C(n4643), .Y(n4641));
   AOI22X1 U5517 ( .A(n2121),  .B(n3843),  .C(n2125),  .D(n3971), .Y(n4643));
   INVX1 U5518 ( .A(w_mem_inst_w_mem[426]), .Y(n3971));
   INVX1 U5519 ( .A(w_mem_inst_w_mem[362]), .Y(n3843));
   NAND2X1 U5520 ( .A(n2119),  .B(n4099), .Y(n4642));
   INVX1 U5521 ( .A(w_mem_inst_w_mem[490]), .Y(n4099));
   NAND3X1 U5522 ( .A(n4644),  .B(n4645),  .C(n4646), .Y(n4640));
   AOI22X1 U5523 ( .A(n4158),  .B(n4035),  .C(n2123),  .D(n3715), .Y(n4646));
   INVX1 U5524 ( .A(w_mem_inst_w_mem[298]), .Y(n3715));
   INVX1 U5525 ( .A(w_mem_inst_w_mem[458]), .Y(n4035));
   NAND2X1 U5526 ( .A(n3106),  .B(n3651), .Y(n4645));
   INVX1 U5527 ( .A(w_mem_inst_w_mem[266]), .Y(n3651));
   AOI22X1 U5528 ( .A(n4160),  .B(n3779),  .C(n4161),  .D(n3907), .Y(n4644));
   INVX1 U5529 ( .A(w_mem_inst_w_mem[394]), .Y(n3907));
   INVX1 U5530 ( .A(w_mem_inst_w_mem[330]), .Y(n3779));
   NAND3X1 U5531 ( .A(n4647),  .B(n4648),  .C(n4649), .Y(n4638));
   AND2X1 U5532 ( .A(n4650),  .B(n4651), .Y(n4649));
   AOI22X1 U5533 ( .A(n4158),  .B(n3523),  .C(n2123),  .D(n3203), .Y(n4651));
   INVX1 U5534 ( .A(w_mem_inst_w_mem[42]), .Y(n3203));
   INVX1 U5535 ( .A(w_mem_inst_w_mem[202]), .Y(n3523));
   AOI22X1 U5536 ( .A(n2121),  .B(n3331),  .C(n2125),  .D(n3459), .Y(n4650));
   INVX1 U5537 ( .A(w_mem_inst_w_mem[170]), .Y(n3459));
   INVX1 U5538 ( .A(w_mem_inst_w_mem[106]), .Y(n3331));
   OAI21X1 U5539 ( .A(n3139),  .B(n2895),  .C(n2117), .Y(n4648));
   INVX1 U5540 ( .A(w_mem_inst_w_mem[10]), .Y(n3139));
   AOI22X1 U5541 ( .A(n2119),  .B(n3587),  .C(n4652),  .D(n4653), .Y(n4647));
   NAND2X1 U5542 ( .A(w_mem_inst_w_mem[138]),  .B(n2894), .Y(n4653));
   AOI21X1 U5543 ( .A(w_mem_inst_w_mem[74]),  .B(n2958),  .C(n4169), .Y(n4652));
   INVX1 U5544 ( .A(w_mem_inst_w_mem[234]), .Y(n3587));
   NAND3X1 U5545 ( .A(n4149),  .B(n4658),  .C(n4659), .Y(n4657));
   AOI22X1 U5546 ( .A(n2121),  .B(n3823),  .C(n2125),  .D(n3951), .Y(n4659));
   INVX1 U5547 ( .A(w_mem_inst_w_mem[416]), .Y(n3951));
   INVX1 U5548 ( .A(w_mem_inst_w_mem[352]), .Y(n3823));
   NAND2X1 U5549 ( .A(n2119),  .B(n4079), .Y(n4658));
   INVX1 U5550 ( .A(w_mem_inst_w_mem[480]), .Y(n4079));
   AND2X1 U5551 ( .A(n4144),  .B(n3111), .Y(n4149));
   INVX1 U5552 ( .A(w_mem_inst_w_ctr_reg[3]), .Y(n3111));
   NAND3X1 U5553 ( .A(n4660),  .B(n4661),  .C(n4662), .Y(n4656));
   AOI22X1 U5554 ( .A(n4158),  .B(n4015),  .C(n2123),  .D(n3695), .Y(n4662));
   INVX1 U5555 ( .A(w_mem_inst_w_mem[288]), .Y(n3695));
   INVX1 U5556 ( .A(w_mem_inst_w_mem[448]), .Y(n4015));
   NAND2X1 U5557 ( .A(n3106),  .B(n3631), .Y(n4661));
   INVX1 U5558 ( .A(w_mem_inst_w_mem[256]), .Y(n3631));
   INVX1 U5559 ( .A(n1953), .Y(n3106));
   AOI22X1 U5560 ( .A(n4160),  .B(n3759),  .C(n4161),  .D(n3887), .Y(n4660));
   INVX1 U5561 ( .A(w_mem_inst_w_mem[384]), .Y(n3887));
   INVX1 U5562 ( .A(n2958), .Y(n4161));
   INVX1 U5563 ( .A(w_mem_inst_w_mem[320]), .Y(n3759));
   INVX1 U5564 ( .A(n2894), .Y(n4160));
   NAND3X1 U5565 ( .A(n4664),  .B(n4665),  .C(n4666), .Y(n4654));
   AND2X1 U5566 ( .A(n4667),  .B(n4668), .Y(n4666));
   AOI22X1 U5567 ( .A(n4158),  .B(n3503),  .C(n2123),  .D(n3183), .Y(n4668));
   INVX1 U5568 ( .A(w_mem_inst_w_mem[32]), .Y(n3183));
   NOR3X1 U5569 ( .A(n3107),  .B(w_mem_inst_w_ctr_reg[0]),  .C(n3109), .Y(n4159));
   INVX1 U5570 ( .A(w_mem_inst_w_mem[192]), .Y(n3503));
   INVX1 U5571 ( .A(n4669), .Y(n4158));
   NAND3X1 U5572 ( .A(n3107),  .B(n3109),  .C(w_mem_inst_w_ctr_reg[0]), .Y(n4669));
   AOI22X1 U5573 ( .A(n2121),  .B(n3311),  .C(n2125),  .D(n3439), .Y(n4667));
   INVX1 U5574 ( .A(w_mem_inst_w_mem[160]), .Y(n3439));
   NOR3X1 U5575 ( .A(w_mem_inst_w_ctr_reg[0]),  .B(w_mem_inst_w_ctr_reg[2]),  .C(n3107), .Y(n4153));
   INVX1 U5576 ( .A(w_mem_inst_w_mem[96]), .Y(n3311));
   NOR3X1 U5577 ( .A(w_mem_inst_w_ctr_reg[0]),  .B(w_mem_inst_w_ctr_reg[1]),  .C(n3109), .Y(n4152));
   OAI21X1 U5578 ( .A(n3118),  .B(n2895),  .C(n2117), .Y(n4665));
   NAND3X1 U5579 ( .A(w_mem_inst_w_ctr_reg[1]),  .B(w_mem_inst_w_ctr_reg[0]),  .C(w_mem_inst_w_ctr_reg[2]), .Y(n4663));
   INVX1 U5580 ( .A(w_mem_inst_w_ctr_reg[4]), .Y(n3113));
   INVX1 U5581 ( .A(w_mem_inst_w_ctr_reg[5]), .Y(n3098));
   INVX1 U5582 ( .A(w_mem_inst_w_mem[0]), .Y(n3118));
   AOI22X1 U5583 ( .A(n2119),  .B(n3567),  .C(n4670),  .D(n4671), .Y(n4664));
   NAND2X1 U5584 ( .A(w_mem_inst_w_mem[128]),  .B(n2894), .Y(n4671));
   AOI21X1 U5585 ( .A(w_mem_inst_w_mem[64]),  .B(n2958),  .C(n4169), .Y(n4670));
   NAND3X1 U5586 ( .A(w_mem_inst_w_ctr_reg[0]),  .B(n3107),  .C(w_mem_inst_w_ctr_reg[2]), .Y(n4445));
   INVX1 U5587 ( .A(w_mem_inst_w_ctr_reg[1]), .Y(n3107));
   NAND3X1 U5588 ( .A(w_mem_inst_w_ctr_reg[0]),  .B(n3109),  .C(w_mem_inst_w_ctr_reg[1]), .Y(n4168));
   INVX1 U5589 ( .A(w_mem_inst_w_ctr_reg[2]), .Y(n3109));
   INVX1 U5590 ( .A(w_mem_inst_w_mem[224]), .Y(n3567));
   NOR3X1 U5591 ( .A(w_mem_inst_w_ctr_reg[1]),  .B(w_mem_inst_w_ctr_reg[2]),  .C(w_mem_inst_w_ctr_reg[0]), .Y(n4154));
   OAI21X1 U5592 ( .A(n4672),  .B(n4673),  .C(n4674), .Y(n6194));
   OAI21X1 U5593 ( .A(a_reg[2]),  .B(b_reg[2]),  .C(c_reg[2]), .Y(n4674));
   INVX1 U5594 ( .A(b_reg[2]), .Y(n4673));
   OAI21X1 U5595 ( .A(n4675),  .B(n4676),  .C(n4677), .Y(n6195));
   OAI21X1 U5596 ( .A(a_reg[9]),  .B(b_reg[9]),  .C(c_reg[9]), .Y(n4677));
   INVX1 U5597 ( .A(b_reg[9]), .Y(n4676));
   INVX1 U5598 ( .A(n4678), .Y(n6196));
   AOI21X1 U5599 ( .A(a_reg[10]),  .B(b_reg[10]),  .C(n4679), .Y(puf_11_wire_3));
   INVX1 U5600 ( .A(n4680), .Y(n4679));
   OAI21X1 U5601 ( .A(a_reg[10]),  .B(b_reg[10]),  .C(c_reg[10]), .Y(n4680));
   OAI21X1 U5602 ( .A(n4681),  .B(n4682),  .C(n4683), .Y(n6197));
   OAI21X1 U5603 ( .A(a_reg[25]),  .B(b_reg[25]),  .C(c_reg[25]), .Y(n4683));
   INVX1 U5604 ( .A(b_reg[25]), .Y(n4682));
   OAI21X1 U5605 ( .A(n4684),  .B(n4685),  .C(n4686), .Y(n6198));
   OAI21X1 U5606 ( .A(a_reg[27]),  .B(b_reg[27]),  .C(c_reg[27]), .Y(n4686));
   INVX1 U5607 ( .A(b_reg[27]), .Y(n4685));
   OAI21X1 U5608 ( .A(n4687),  .B(n4688),  .C(n4689), .Y(n6199));
   OAI21X1 U5609 ( .A(a_reg[29]),  .B(b_reg[29]),  .C(c_reg[29]), .Y(n4689));
   INVX1 U5610 ( .A(b_reg[29]), .Y(n4688));
   NAND2X1 U5611 ( .A(n3049),  .B(n4690), .Y(n1755));
   NAND3X1 U5612 ( .A(n4691),  .B(n3100),  .C(sha256_ctrl_reg[0]), .Y(n4690));
   NAND3X1 U5613 ( .A(n6068),  .B(n4692),  .C(t_ctr_reg[3]), .Y(n4691));
   AOI21X1 U5614 ( .A(n4693),  .B(n4694),  .C(n4695), .Y(n1754));
   NAND3X1 U5615 ( .A(n6068),  .B(n2980),  .C(t_ctr_reg[3]), .Y(n4694));
   NAND2X1 U5616 ( .A(sha256_ctrl_reg[1]),  .B(n3100), .Y(n4693));
   NAND2X1 U5617 ( .A(n2887),  .B(n4697), .Y(n1753));
   NAND3X1 U5618 ( .A(n4698),  .B(n3100),  .C(digest_valid), .Y(n4697));
   OAI21X1 U5619 ( .A(next),  .B(init),  .C(n4695), .Y(n4698));
   MUX2X1 U5620 ( .A(n2102),  .B(n2126),  .S(n4700), .Y(n1752));
   OAI21X1 U5621 ( .A(n4701),  .B(n2126),  .C(n4702), .Y(n1751));
   NAND2X1 U5622 ( .A(N1615),  .B(n2979), .Y(n4702));
   OAI21X1 U5623 ( .A(n4703),  .B(n2126),  .C(n4704), .Y(n1750));
   NAND2X1 U5624 ( .A(N1616),  .B(n2980), .Y(n4704));
   OAI21X1 U5625 ( .A(n4705),  .B(n2126),  .C(n4706), .Y(n1749));
   NAND2X1 U5626 ( .A(N1617),  .B(n2980), .Y(n4706));
   OAI21X1 U5627 ( .A(n4707),  .B(n2126),  .C(n4708), .Y(n1748));
   NAND2X1 U5628 ( .A(N1618),  .B(n2980), .Y(n4708));
   MUX2X1 U5629 ( .A(n4710),  .B(n4709),  .S(n4711), .Y(n1747));
   NAND2X1 U5630 ( .A(add_420_carry[5]),  .B(n2977), .Y(n4710));
   INVX1 U5631 ( .A(n4712), .Y(n4709));
   OAI21X1 U5632 ( .A(n2102),  .B(add_420_carry[5]),  .C(n2126), .Y(n4712));
   OAI21X1 U5633 ( .A(n3083),  .B(n4714),  .C(n2264), .Y(n1746));
   INVX1 U5634 ( .A(digest[128]), .Y(n4714));
   NAND2X1 U5635 ( .A(n4716),  .B(n4717), .Y(n1745));
   NAND2X1 U5636 ( .A(d_reg[0]),  .B(n3089), .Y(n4717));
   AOI22X1 U5637 ( .A(c_reg[0]),  .B(n2977),  .C(n4718),  .D(digest[128]), .Y(n4716));
   NAND3X1 U5638 ( .A(n4719),  .B(n3090),  .C(n4720), .Y(n1744));
   AOI22X1 U5639 ( .A(c_reg[1]),  .B(n2977),  .C(d_reg[1]),  .D(n3088), .Y(n4720));
   NAND2X1 U5640 ( .A(digest[129]),  .B(n3050), .Y(n4719));
   NAND2X1 U5641 ( .A(n4721),  .B(n4722), .Y(n1743));
   NAND2X1 U5642 ( .A(d_reg[2]),  .B(n3089), .Y(n4722));
   AOI22X1 U5643 ( .A(c_reg[2]),  .B(n2978),  .C(digest[130]),  .D(n4718), .Y(n4721));
   NAND3X1 U5644 ( .A(n4723),  .B(n3091),  .C(n4724), .Y(n1742));
   AOI22X1 U5645 ( .A(c_reg[3]),  .B(n2980),  .C(d_reg[3]),  .D(n3089), .Y(n4724));
   NAND2X1 U5646 ( .A(digest[131]),  .B(n3050), .Y(n4723));
   NAND3X1 U5647 ( .A(n4725),  .B(n3091),  .C(n4726), .Y(n1741));
   AOI22X1 U5648 ( .A(c_reg[4]),  .B(n2977),  .C(d_reg[4]),  .D(n3089), .Y(n4726));
   NAND2X1 U5649 ( .A(digest[132]),  .B(n3050), .Y(n4725));
   NAND3X1 U5650 ( .A(n4727),  .B(n3090),  .C(n4728), .Y(n1740));
   AOI22X1 U5651 ( .A(c_reg[5]),  .B(n2979),  .C(d_reg[5]),  .D(n3089), .Y(n4728));
   NAND2X1 U5652 ( .A(digest[133]),  .B(n3050), .Y(n4727));
   NAND2X1 U5653 ( .A(n4729),  .B(n4730), .Y(n1739));
   NAND2X1 U5654 ( .A(d_reg[6]),  .B(n3088), .Y(n4730));
   AOI22X1 U5655 ( .A(c_reg[6]),  .B(n2979),  .C(digest[134]),  .D(n4718), .Y(n4729));
   NAND2X1 U5656 ( .A(n4731),  .B(n4732), .Y(n1738));
   NAND2X1 U5657 ( .A(d_reg[7]),  .B(n3089), .Y(n4732));
   AOI22X1 U5658 ( .A(c_reg[7]),  .B(n2978),  .C(digest[135]),  .D(n4718), .Y(n4731));
   NAND3X1 U5659 ( .A(n4733),  .B(n3091),  .C(n4734), .Y(n1737));
   AOI22X1 U5660 ( .A(c_reg[8]),  .B(n2978),  .C(d_reg[8]),  .D(n3089), .Y(n4734));
   NAND2X1 U5661 ( .A(digest[136]),  .B(n3050), .Y(n4733));
   NAND2X1 U5662 ( .A(n4735),  .B(n4736), .Y(n1736));
   NAND2X1 U5663 ( .A(d_reg[9]),  .B(n3089), .Y(n4736));
   AOI22X1 U5664 ( .A(c_reg[9]),  .B(n2978),  .C(digest[137]),  .D(n4718), .Y(n4735));
   NAND3X1 U5665 ( .A(n4737),  .B(n3091),  .C(n4738), .Y(n1735));
   AOI22X1 U5666 ( .A(c_reg[10]),  .B(n2978),  .C(d_reg[10]),  .D(n3089), .Y(n4738));
   NAND2X1 U5667 ( .A(digest[138]),  .B(n3050), .Y(n4737));
   NAND2X1 U5668 ( .A(n4739),  .B(n4740), .Y(n1734));
   NAND2X1 U5669 ( .A(d_reg[11]),  .B(n3089), .Y(n4740));
   AOI22X1 U5670 ( .A(c_reg[11]),  .B(n2980),  .C(digest[139]),  .D(n4718), .Y(n4739));
   NAND3X1 U5671 ( .A(n4741),  .B(n3091),  .C(n4742), .Y(n1733));
   AOI22X1 U5672 ( .A(c_reg[12]),  .B(n2979),  .C(d_reg[12]),  .D(n3089), .Y(n4742));
   NAND2X1 U5673 ( .A(digest[140]),  .B(n3050), .Y(n4741));
   NAND3X1 U5674 ( .A(n4743),  .B(n3091),  .C(n4744), .Y(n1732));
   AOI22X1 U5675 ( .A(c_reg[13]),  .B(n2977),  .C(d_reg[13]),  .D(n3089), .Y(n4744));
   NAND2X1 U5676 ( .A(digest[141]),  .B(n3050), .Y(n4743));
   NAND3X1 U5677 ( .A(n4745),  .B(n3091),  .C(n4746), .Y(n1731));
   AOI22X1 U5678 ( .A(c_reg[14]),  .B(n2979),  .C(d_reg[14]),  .D(n3089), .Y(n4746));
   NAND2X1 U5679 ( .A(digest[142]),  .B(n3050), .Y(n4745));
   NAND3X1 U5680 ( .A(n4747),  .B(n3091),  .C(n4748), .Y(n1730));
   AOI22X1 U5681 ( .A(c_reg[15]),  .B(n2978),  .C(d_reg[15]),  .D(n3089), .Y(n4748));
   NAND2X1 U5682 ( .A(digest[143]),  .B(n3050), .Y(n4747));
   NAND3X1 U5683 ( .A(n4749),  .B(n3091),  .C(n4750), .Y(n1729));
   AOI22X1 U5684 ( .A(c_reg[16]),  .B(n2980),  .C(d_reg[16]),  .D(n3089), .Y(n4750));
   NAND2X1 U5685 ( .A(digest[144]),  .B(n3048), .Y(n4749));
   NAND3X1 U5686 ( .A(n4751),  .B(n3091),  .C(n4752), .Y(n1728));
   AOI22X1 U5687 ( .A(c_reg[17]),  .B(n2979),  .C(d_reg[17]),  .D(n3088), .Y(n4752));
   NAND2X1 U5688 ( .A(digest[145]),  .B(n3048), .Y(n4751));
   NAND3X1 U5689 ( .A(n4753),  .B(n3091),  .C(n4754), .Y(n1727));
   AOI22X1 U5690 ( .A(c_reg[18]),  .B(n2977),  .C(d_reg[18]),  .D(n3089), .Y(n4754));
   NAND2X1 U5691 ( .A(digest[146]),  .B(n3048), .Y(n4753));
   NAND3X1 U5692 ( .A(n4755),  .B(n3091),  .C(n4756), .Y(n1726));
   AOI22X1 U5693 ( .A(c_reg[19]),  .B(n2977),  .C(d_reg[19]),  .D(n3088), .Y(n4756));
   NAND2X1 U5694 ( .A(digest[147]),  .B(n3048), .Y(n4755));
   NAND2X1 U5695 ( .A(n4757),  .B(n4758), .Y(n1725));
   NAND2X1 U5696 ( .A(d_reg[20]),  .B(n3089), .Y(n4758));
   AOI22X1 U5697 ( .A(c_reg[20]),  .B(n2978),  .C(digest[148]),  .D(n4718), .Y(n4757));
   NAND2X1 U5698 ( .A(n4759),  .B(n4760), .Y(n1724));
   NAND2X1 U5699 ( .A(d_reg[21]),  .B(n3088), .Y(n4760));
   AOI22X1 U5700 ( .A(c_reg[21]),  .B(n2980),  .C(digest[149]),  .D(n4718), .Y(n4759));
   NAND3X1 U5701 ( .A(n4761),  .B(n3091),  .C(n4762), .Y(n1723));
   AOI22X1 U5702 ( .A(c_reg[22]),  .B(n2979),  .C(d_reg[22]),  .D(n3088), .Y(n4762));
   NAND2X1 U5703 ( .A(digest[150]),  .B(n3048), .Y(n4761));
   NAND2X1 U5704 ( .A(n4763),  .B(n4764), .Y(n1722));
   NAND2X1 U5705 ( .A(d_reg[23]),  .B(n3088), .Y(n4764));
   AOI22X1 U5706 ( .A(c_reg[23]),  .B(n2977),  .C(digest[151]),  .D(n4718), .Y(n4763));
   NAND3X1 U5707 ( .A(n4765),  .B(n3091),  .C(n4766), .Y(n1721));
   AOI22X1 U5708 ( .A(c_reg[24]),  .B(n2980),  .C(d_reg[24]),  .D(n3088), .Y(n4766));
   NAND2X1 U5709 ( .A(digest[152]),  .B(n3048), .Y(n4765));
   NAND2X1 U5710 ( .A(n4767),  .B(n4768), .Y(n1720));
   NAND2X1 U5711 ( .A(d_reg[25]),  .B(n3089), .Y(n4768));
   AOI22X1 U5712 ( .A(c_reg[25]),  .B(n2980),  .C(digest[153]),  .D(n4718), .Y(n4767));
   NAND3X1 U5713 ( .A(n4769),  .B(n3091),  .C(n4770), .Y(n1719));
   AOI22X1 U5714 ( .A(c_reg[26]),  .B(n2980),  .C(d_reg[26]),  .D(n3088), .Y(n4770));
   NAND2X1 U5715 ( .A(digest[154]),  .B(n3048), .Y(n4769));
   NAND2X1 U5716 ( .A(n4771),  .B(n4772), .Y(n1718));
   NAND2X1 U5717 ( .A(d_reg[27]),  .B(n3089), .Y(n4772));
   AOI22X1 U5718 ( .A(c_reg[27]),  .B(n2979),  .C(digest[155]),  .D(n4718), .Y(n4771));
   NAND2X1 U5719 ( .A(n4773),  .B(n4774), .Y(n1717));
   NAND2X1 U5720 ( .A(d_reg[28]),  .B(n3089), .Y(n4774));
   AOI22X1 U5721 ( .A(c_reg[28]),  .B(n2977),  .C(digest[156]),  .D(n4718), .Y(n4773));
   NAND3X1 U5722 ( .A(n4775),  .B(n3091),  .C(n4776), .Y(n1716));
   AOI22X1 U5723 ( .A(c_reg[29]),  .B(n2980),  .C(d_reg[29]),  .D(n3088), .Y(n4776));
   NAND2X1 U5724 ( .A(digest[157]),  .B(n3048), .Y(n4775));
   NAND2X1 U5725 ( .A(n4777),  .B(n4778), .Y(n1715));
   NAND2X1 U5726 ( .A(d_reg[30]),  .B(n3089), .Y(n4778));
   AOI22X1 U5727 ( .A(c_reg[30]),  .B(n2978),  .C(digest[158]),  .D(n4718), .Y(n4777));
   NAND3X1 U5728 ( .A(n4779),  .B(n3091),  .C(n4780), .Y(n1714));
   AOI22X1 U5729 ( .A(c_reg[31]),  .B(n2979),  .C(d_reg[31]),  .D(n3088), .Y(n4780));
   NAND2X1 U5730 ( .A(digest[159]),  .B(n3048), .Y(n4779));
   OAI21X1 U5731 ( .A(n3082),  .B(n4781),  .C(n2647), .Y(n1713));
   AOI21X1 U5732 ( .A(N647),  .B(n3085),  .C(n4783), .Y(n4782));
   INVX1 U5733 ( .A(digest[129]), .Y(n4781));
   OAI21X1 U5734 ( .A(n3083),  .B(n4784),  .C(n2198), .Y(n1712));
   INVX1 U5735 ( .A(digest[130]), .Y(n4784));
   OAI21X1 U5736 ( .A(n4713),  .B(n4786),  .C(n2532), .Y(n1711));
   AOI21X1 U5737 ( .A(N649),  .B(n3085),  .C(n4783), .Y(n4787));
   INVX1 U5738 ( .A(digest[131]), .Y(n4786));
   OAI21X1 U5739 ( .A(n3082),  .B(n4788),  .C(n2710), .Y(n1710));
   AOI21X1 U5740 ( .A(N650),  .B(n3086),  .C(n4783), .Y(n4789));
   INVX1 U5741 ( .A(digest[132]), .Y(n4788));
   OAI21X1 U5742 ( .A(n3082),  .B(n4790),  .C(n2774), .Y(n1709));
   AOI21X1 U5743 ( .A(N651),  .B(n3085),  .C(n4783), .Y(n4791));
   INVX1 U5744 ( .A(digest[133]), .Y(n4790));
   OAI21X1 U5745 ( .A(n4713),  .B(n4792),  .C(n2228), .Y(n1708));
   INVX1 U5746 ( .A(digest[134]), .Y(n4792));
   OAI21X1 U5747 ( .A(n3082),  .B(n4794),  .C(n2375), .Y(n1707));
   INVX1 U5748 ( .A(digest[135]), .Y(n4794));
   OAI21X1 U5749 ( .A(n4713),  .B(n4796),  .C(n2837), .Y(n1706));
   AOI21X1 U5750 ( .A(N654),  .B(n3086),  .C(n4783), .Y(n4797));
   INVX1 U5751 ( .A(digest[136]), .Y(n4796));
   OAI21X1 U5752 ( .A(n4713),  .B(n4798),  .C(n2663), .Y(n1705));
   INVX1 U5753 ( .A(digest[137]), .Y(n4798));
   OAI21X1 U5754 ( .A(n3082),  .B(n4800),  .C(n2944), .Y(n1704));
   AOI21X1 U5755 ( .A(N656),  .B(n3087),  .C(n4783), .Y(n4801));
   INVX1 U5756 ( .A(digest[138]), .Y(n4800));
   OAI21X1 U5757 ( .A(n3083),  .B(n4802),  .C(n2726), .Y(n1703));
   INVX1 U5758 ( .A(digest[139]), .Y(n4802));
   OAI21X1 U5759 ( .A(n4713),  .B(n4804),  .C(n2263), .Y(n1702));
   AOI21X1 U5760 ( .A(N658),  .B(n3086),  .C(n3093), .Y(n4805));
   INVX1 U5761 ( .A(digest[140]), .Y(n4804));
   OAI21X1 U5762 ( .A(n3083),  .B(n4806),  .C(n2314), .Y(n1701));
   AOI21X1 U5763 ( .A(N659),  .B(n3087),  .C(n3093), .Y(n4807));
   INVX1 U5764 ( .A(digest[141]), .Y(n4806));
   OAI21X1 U5765 ( .A(n3083),  .B(n4808),  .C(n2368), .Y(n1700));
   AOI21X1 U5766 ( .A(N660),  .B(n3086),  .C(n3093), .Y(n4809));
   INVX1 U5767 ( .A(digest[142]), .Y(n4808));
   OAI21X1 U5768 ( .A(n4713),  .B(n4810),  .C(n2423), .Y(n1699));
   AOI21X1 U5769 ( .A(N661),  .B(n3085),  .C(n3093), .Y(n4811));
   INVX1 U5770 ( .A(digest[143]), .Y(n4810));
   OAI21X1 U5771 ( .A(n3082),  .B(n4812),  .C(n2478), .Y(n1698));
   AOI21X1 U5772 ( .A(N662),  .B(n3085),  .C(n3093), .Y(n4813));
   INVX1 U5773 ( .A(digest[144]), .Y(n4812));
   OAI21X1 U5774 ( .A(n4713),  .B(n4814),  .C(n2533), .Y(n1697));
   AOI21X1 U5775 ( .A(N663),  .B(n3086),  .C(n3093), .Y(n4815));
   INVX1 U5776 ( .A(digest[145]), .Y(n4814));
   OAI21X1 U5777 ( .A(n3082),  .B(n4816),  .C(n2590), .Y(n1696));
   AOI21X1 U5778 ( .A(N664),  .B(n3087),  .C(n3093), .Y(n4817));
   INVX1 U5779 ( .A(digest[146]), .Y(n4816));
   OAI21X1 U5780 ( .A(n4713),  .B(n4818),  .C(n2648), .Y(n1695));
   AOI21X1 U5781 ( .A(N665),  .B(n3086),  .C(n3093), .Y(n4819));
   INVX1 U5782 ( .A(digest[147]), .Y(n4818));
   OAI21X1 U5783 ( .A(n3083),  .B(n4820),  .C(n2790), .Y(n1694));
   INVX1 U5784 ( .A(digest[148]), .Y(n4820));
   OAI21X1 U5785 ( .A(n3083),  .B(n4822),  .C(n2321), .Y(n1693));
   INVX1 U5786 ( .A(digest[149]), .Y(n4822));
   OAI21X1 U5787 ( .A(n4713),  .B(n4824),  .C(n2711), .Y(n1692));
   AOI21X1 U5788 ( .A(N668),  .B(n3086),  .C(n3093), .Y(n4825));
   INVX1 U5789 ( .A(digest[150]), .Y(n4824));
   OAI21X1 U5790 ( .A(n3083),  .B(n4826),  .C(n2376), .Y(n1691));
   INVX1 U5791 ( .A(digest[151]), .Y(n4826));
   OAI21X1 U5792 ( .A(n3082),  .B(n4828),  .C(n2775), .Y(n1690));
   AOI21X1 U5793 ( .A(N670),  .B(n3085),  .C(n3093), .Y(n4829));
   INVX1 U5794 ( .A(digest[152]), .Y(n4828));
   OAI21X1 U5795 ( .A(n4713),  .B(n4830),  .C(n2432), .Y(n1689));
   INVX1 U5796 ( .A(digest[153]), .Y(n4830));
   OAI21X1 U5797 ( .A(n3082),  .B(n4832),  .C(n2838), .Y(n1688));
   AOI21X1 U5798 ( .A(N672),  .B(n3086),  .C(n3093), .Y(n4833));
   INVX1 U5799 ( .A(digest[154]), .Y(n4832));
   OAI21X1 U5800 ( .A(n4713),  .B(n4834),  .C(n2488), .Y(n1687));
   INVX1 U5801 ( .A(digest[155]), .Y(n4834));
   OAI21X1 U5802 ( .A(n3082),  .B(n4836),  .C(n2601), .Y(n1686));
   INVX1 U5803 ( .A(digest[156]), .Y(n4836));
   OAI21X1 U5804 ( .A(n4713),  .B(n4838),  .C(n2945), .Y(n1685));
   AOI21X1 U5805 ( .A(N675),  .B(n3086),  .C(n3093), .Y(n4839));
   INVX1 U5806 ( .A(digest[157]), .Y(n4838));
   OAI21X1 U5807 ( .A(n4713),  .B(n4840),  .C(n2546), .Y(n1684));
   INVX1 U5808 ( .A(digest[158]), .Y(n4840));
   OAI21X1 U5809 ( .A(n3082),  .B(n4842),  .C(n4843), .Y(n1683));
   AOI21X1 U5810 ( .A(N677),  .B(n3087),  .C(n3093), .Y(n4843));
   INVX1 U5811 ( .A(digest[159]), .Y(n4842));
   NAND3X1 U5812 ( .A(n4844),  .B(n3090),  .C(n4845), .Y(n1682));
   AOI22X1 U5813 ( .A(N1579),  .B(n2978),  .C(e_reg[0]),  .D(n3088), .Y(n4845));
   NAND2X1 U5814 ( .A(digest[96]),  .B(n3048), .Y(n4844));
   NAND3X1 U5815 ( .A(n4846),  .B(n3090),  .C(n4847), .Y(n1681));
   AOI22X1 U5816 ( .A(N1580),  .B(n2980),  .C(e_reg[1]),  .D(n3089), .Y(n4847));
   NAND2X1 U5817 ( .A(digest[97]),  .B(n3048), .Y(n4846));
   NAND3X1 U5818 ( .A(n4848),  .B(n3090),  .C(n4849), .Y(n1680));
   AOI22X1 U5819 ( .A(N1581),  .B(n2979),  .C(e_reg[2]),  .D(n3088), .Y(n4849));
   NAND2X1 U5820 ( .A(digest[98]),  .B(n3048), .Y(n4848));
   NAND3X1 U5821 ( .A(n4850),  .B(n3090),  .C(n4851), .Y(n1679));
   AOI22X1 U5822 ( .A(N1582),  .B(n2977),  .C(e_reg[3]),  .D(n3088), .Y(n4851));
   NAND2X1 U5823 ( .A(digest[99]),  .B(n3048), .Y(n4850));
   NAND3X1 U5824 ( .A(n4852),  .B(n3090),  .C(n4853), .Y(n1678));
   AOI22X1 U5825 ( .A(N1583),  .B(n2979),  .C(e_reg[4]),  .D(n3088), .Y(n4853));
   NAND2X1 U5826 ( .A(digest[100]),  .B(n3048), .Y(n4852));
   NAND3X1 U5827 ( .A(n4854),  .B(n3090),  .C(n4855), .Y(n1677));
   AOI22X1 U5828 ( .A(N1584),  .B(n2979),  .C(e_reg[5]),  .D(n3089), .Y(n4855));
   NAND2X1 U5829 ( .A(digest[101]),  .B(n3048), .Y(n4854));
   NAND3X1 U5830 ( .A(n4856),  .B(n3090),  .C(n4857), .Y(n1676));
   AOI22X1 U5831 ( .A(N1585),  .B(n2979),  .C(e_reg[6]),  .D(n3089), .Y(n4857));
   NAND2X1 U5832 ( .A(digest[102]),  .B(n3048), .Y(n4856));
   OAI21X1 U5833 ( .A(n2126),  .B(n4858),  .C(n4859), .Y(n1675));
   AOI22X1 U5834 ( .A(N1586),  .B(n2979),  .C(digest[103]),  .D(n4718), .Y(n4859));
   OAI21X1 U5835 ( .A(n2126),  .B(n4860),  .C(n4861), .Y(n1674));
   AOI22X1 U5836 ( .A(N1587),  .B(n2979),  .C(digest[104]),  .D(n4718), .Y(n4861));
   NAND3X1 U5837 ( .A(n4862),  .B(n3090),  .C(n4863), .Y(n1673));
   AOI22X1 U5838 ( .A(N1588),  .B(n2979),  .C(e_reg[9]),  .D(n3089), .Y(n4863));
   NAND2X1 U5839 ( .A(digest[105]),  .B(n3048), .Y(n4862));
   OAI21X1 U5840 ( .A(n2126),  .B(n4864),  .C(n4865), .Y(n1672));
   AOI22X1 U5841 ( .A(N1589),  .B(n2979),  .C(digest[106]),  .D(n4718), .Y(n4865));
   OAI21X1 U5842 ( .A(n2126),  .B(n4866),  .C(n4867), .Y(n1671));
   AOI22X1 U5843 ( .A(N1590),  .B(n2979),  .C(digest[107]),  .D(n4718), .Y(n4867));
   NAND3X1 U5844 ( .A(n4868),  .B(n3090),  .C(n4869), .Y(n1670));
   AOI22X1 U5845 ( .A(N1591),  .B(n2979),  .C(e_reg[12]),  .D(n3088), .Y(n4869));
   NAND2X1 U5846 ( .A(digest[108]),  .B(n3046), .Y(n4868));
   OAI21X1 U5847 ( .A(n2126),  .B(n4870),  .C(n4871), .Y(n1669));
   AOI22X1 U5848 ( .A(N1592),  .B(n2979),  .C(digest[109]),  .D(n4718), .Y(n4871));
   NAND3X1 U5849 ( .A(n4872),  .B(n3090),  .C(n4873), .Y(n1668));
   AOI22X1 U5850 ( .A(N1593),  .B(n2979),  .C(e_reg[14]),  .D(n3088), .Y(n4873));
   NAND2X1 U5851 ( .A(digest[110]),  .B(n3050), .Y(n4872));
   OAI21X1 U5852 ( .A(n2126),  .B(n4874),  .C(n4875), .Y(n1667));
   AOI22X1 U5853 ( .A(N1594),  .B(n2979),  .C(digest[111]),  .D(n4718), .Y(n4875));
   OAI21X1 U5854 ( .A(n2126),  .B(n4876),  .C(n4877), .Y(n1666));
   AOI22X1 U5855 ( .A(N1595),  .B(n2979),  .C(digest[112]),  .D(n4718), .Y(n4877));
   NAND3X1 U5856 ( .A(n4878),  .B(n3090),  .C(n4879), .Y(n1665));
   AOI22X1 U5857 ( .A(N1596),  .B(n2979),  .C(e_reg[17]),  .D(n3088), .Y(n4879));
   NAND2X1 U5858 ( .A(digest[113]),  .B(n3041), .Y(n4878));
   NAND3X1 U5859 ( .A(n4880),  .B(n3090),  .C(n4881), .Y(n1664));
   AOI22X1 U5860 ( .A(N1597),  .B(n2978),  .C(e_reg[18]),  .D(n3089), .Y(n4881));
   NAND2X1 U5861 ( .A(digest[114]),  .B(n3048), .Y(n4880));
   NAND3X1 U5862 ( .A(n4882),  .B(n3090),  .C(n4883), .Y(n1663));
   AOI22X1 U5863 ( .A(N1598),  .B(n2978),  .C(e_reg[19]),  .D(n3088), .Y(n4883));
   NAND2X1 U5864 ( .A(digest[115]),  .B(n3039), .Y(n4882));
   OAI21X1 U5865 ( .A(n2126),  .B(n4884),  .C(n4885), .Y(n1662));
   AOI22X1 U5866 ( .A(N1599),  .B(n2978),  .C(digest[116]),  .D(n4718), .Y(n4885));
   OAI21X1 U5867 ( .A(n2126),  .B(n4886),  .C(n4887), .Y(n1661));
   AOI22X1 U5868 ( .A(N1600),  .B(n2978),  .C(digest[117]),  .D(n4718), .Y(n4887));
   OAI21X1 U5869 ( .A(n2126),  .B(n4888),  .C(n4889), .Y(n1660));
   AOI22X1 U5870 ( .A(N1601),  .B(n2978),  .C(digest[118]),  .D(n4718), .Y(n4889));
   OAI21X1 U5871 ( .A(n2126),  .B(n4890),  .C(n4891), .Y(n1659));
   AOI22X1 U5872 ( .A(N1602),  .B(n2978),  .C(digest[119]),  .D(n4718), .Y(n4891));
   NAND3X1 U5873 ( .A(n4892),  .B(n3090),  .C(n4893), .Y(n1658));
   AOI22X1 U5874 ( .A(N1603),  .B(n2978),  .C(e_reg[24]),  .D(n3088), .Y(n4893));
   NAND2X1 U5875 ( .A(digest[120]),  .B(n3037), .Y(n4892));
   OAI21X1 U5876 ( .A(n2126),  .B(n4894),  .C(n4895), .Y(n1657));
   AOI22X1 U5877 ( .A(N1604),  .B(n2979),  .C(digest[121]),  .D(n4718), .Y(n4895));
   OAI21X1 U5878 ( .A(n2126),  .B(n4896),  .C(n4897), .Y(n1656));
   AOI22X1 U5879 ( .A(N1605),  .B(n2978),  .C(digest[122]),  .D(n4718), .Y(n4897));
   OAI21X1 U5880 ( .A(n2126),  .B(n4898),  .C(n4899), .Y(n1655));
   AOI22X1 U5881 ( .A(N1606),  .B(n2978),  .C(digest[123]),  .D(n4718), .Y(n4899));
   NAND3X1 U5882 ( .A(n4900),  .B(n3091),  .C(n4901), .Y(n1654));
   AOI22X1 U5883 ( .A(N1607),  .B(n2978),  .C(e_reg[28]),  .D(n3088), .Y(n4901));
   NAND2X1 U5884 ( .A(digest[124]),  .B(n3018), .Y(n4900));
   OAI21X1 U5885 ( .A(n2126),  .B(n4902),  .C(n4903), .Y(n1653));
   AOI22X1 U5886 ( .A(N1608),  .B(n2978),  .C(digest[125]),  .D(n4718), .Y(n4903));
   NAND3X1 U5887 ( .A(n4904),  .B(n3090),  .C(n4905), .Y(n1652));
   AOI22X1 U5888 ( .A(N1609),  .B(n2978),  .C(e_reg[30]),  .D(n3089), .Y(n4905));
   NAND2X1 U5889 ( .A(digest[126]),  .B(n3034), .Y(n4904));
   OAI21X1 U5890 ( .A(n2126),  .B(n4906),  .C(n4907), .Y(n1651));
   AOI22X1 U5891 ( .A(N1610),  .B(n2978),  .C(digest[127]),  .D(n4718), .Y(n4907));
   OAI21X1 U5892 ( .A(n3082),  .B(n4908),  .C(n4909), .Y(n1650));
   AOI21X1 U5893 ( .A(N678),  .B(n3087),  .C(n3093), .Y(n4909));
   INVX1 U5894 ( .A(digest[96]), .Y(n4908));
   OAI21X1 U5895 ( .A(n4713),  .B(n4910),  .C(n2168), .Y(n1649));
   AOI21X1 U5896 ( .A(N679),  .B(n3086),  .C(n4783), .Y(n4911));
   INVX1 U5897 ( .A(digest[97]), .Y(n4910));
   OAI21X1 U5898 ( .A(n4713),  .B(n4912),  .C(n2189), .Y(n1648));
   AOI21X1 U5899 ( .A(N680),  .B(n3085),  .C(n4783), .Y(n4913));
   INVX1 U5900 ( .A(digest[98]), .Y(n4912));
   OAI21X1 U5901 ( .A(n3082),  .B(n4914),  .C(n2305), .Y(n1647));
   AOI21X1 U5902 ( .A(N681),  .B(n3087),  .C(n3093), .Y(n4915));
   INVX1 U5903 ( .A(digest[99]), .Y(n4914));
   OAI21X1 U5904 ( .A(n3082),  .B(n4916),  .C(n2359), .Y(n1646));
   AOI21X1 U5905 ( .A(N682),  .B(n3085),  .C(n4783), .Y(n4917));
   INVX1 U5906 ( .A(digest[100]), .Y(n4916));
   OAI21X1 U5907 ( .A(n3083),  .B(n4918),  .C(n2415), .Y(n1645));
   AOI21X1 U5908 ( .A(N683),  .B(n3086),  .C(n4783), .Y(n4919));
   INVX1 U5909 ( .A(digest[101]), .Y(n4918));
   OAI21X1 U5910 ( .A(n3083),  .B(n4920),  .C(n2524), .Y(n1644));
   AOI21X1 U5911 ( .A(N684),  .B(n3085),  .C(n4783), .Y(n4921));
   INVX1 U5912 ( .A(digest[102]), .Y(n4920));
   OAI21X1 U5913 ( .A(n3082),  .B(n4922),  .C(n4923), .Y(n1643));
   NAND2X1 U5914 ( .A(N685),  .B(n3087), .Y(n4923));
   INVX1 U5915 ( .A(digest[103]), .Y(n4922));
   OAI21X1 U5916 ( .A(n4713),  .B(n4924),  .C(n2128), .Y(n1642));
   INVX1 U5917 ( .A(digest[104]), .Y(n4924));
   OAI21X1 U5918 ( .A(n4713),  .B(n4926),  .C(n2582), .Y(n1641));
   AOI21X1 U5919 ( .A(N687),  .B(n3085),  .C(n3093), .Y(n4927));
   INVX1 U5920 ( .A(digest[105]), .Y(n4926));
   OAI21X1 U5921 ( .A(n3083),  .B(n4928),  .C(n2138), .Y(n1640));
   INVX1 U5922 ( .A(digest[106]), .Y(n4928));
   OAI21X1 U5923 ( .A(n3082),  .B(n4930),  .C(n2721), .Y(n1639));
   INVX1 U5924 ( .A(digest[107]), .Y(n4930));
   OAI21X1 U5925 ( .A(n3082),  .B(n4932),  .C(n2215), .Y(n1638));
   AOI21X1 U5926 ( .A(N690),  .B(n3085),  .C(n3093), .Y(n4933));
   INVX1 U5927 ( .A(digest[108]), .Y(n4932));
   OAI21X1 U5928 ( .A(n3083),  .B(n4934),  .C(n4935), .Y(n1637));
   NAND2X1 U5929 ( .A(N691),  .B(n3085), .Y(n4935));
   INVX1 U5930 ( .A(digest[109]), .Y(n4934));
   OAI21X1 U5931 ( .A(n3083),  .B(n4936),  .C(n2257), .Y(n1636));
   AOI21X1 U5932 ( .A(N692),  .B(n3087),  .C(n3093), .Y(n4937));
   INVX1 U5933 ( .A(digest[110]), .Y(n4936));
   OAI21X1 U5934 ( .A(n3083),  .B(n4938),  .C(n2151), .Y(n1635));
   INVX1 U5935 ( .A(digest[111]), .Y(n4938));
   OAI21X1 U5936 ( .A(n3083),  .B(n4940),  .C(n2896), .Y(n1634));
   INVX1 U5937 ( .A(digest[112]), .Y(n4940));
   OAI21X1 U5938 ( .A(n3083),  .B(n4942),  .C(n2639), .Y(n1633));
   AOI21X1 U5939 ( .A(N695),  .B(n3085),  .C(n3093), .Y(n4943));
   INVX1 U5940 ( .A(digest[113]), .Y(n4942));
   OAI21X1 U5941 ( .A(n3083),  .B(n4944),  .C(n2765), .Y(n1632));
   AOI21X1 U5942 ( .A(N696),  .B(n3085),  .C(n4783), .Y(n4945));
   INVX1 U5943 ( .A(digest[114]), .Y(n4944));
   OAI21X1 U5944 ( .A(n3083),  .B(n4946),  .C(n2828), .Y(n1631));
   AOI21X1 U5945 ( .A(N697),  .B(n3086),  .C(n3093), .Y(n4947));
   INVX1 U5946 ( .A(digest[115]), .Y(n4946));
   OAI21X1 U5947 ( .A(n3083),  .B(n4948),  .C(n2129), .Y(n1630));
   INVX1 U5948 ( .A(digest[116]), .Y(n4948));
   OAI21X1 U5949 ( .A(n3083),  .B(n4950),  .C(n2139), .Y(n1629));
   INVX1 U5950 ( .A(digest[117]), .Y(n4950));
   OAI21X1 U5951 ( .A(n3083),  .B(n4952),  .C(n2171), .Y(n1628));
   INVX1 U5952 ( .A(digest[118]), .Y(n4952));
   OAI21X1 U5953 ( .A(n3083),  .B(n4954),  .C(n2193), .Y(n1627));
   INVX1 U5954 ( .A(digest[119]), .Y(n4954));
   OAI21X1 U5955 ( .A(n3083),  .B(n4956),  .C(n2306), .Y(n1626));
   AOI21X1 U5956 ( .A(N702),  .B(n3086),  .C(n3093), .Y(n4957));
   INVX1 U5957 ( .A(digest[120]), .Y(n4956));
   OAI21X1 U5958 ( .A(n3082),  .B(n4958),  .C(n2152), .Y(n1625));
   INVX1 U5959 ( .A(digest[121]), .Y(n4958));
   OAI21X1 U5960 ( .A(n3083),  .B(n4960),  .C(n2221), .Y(n1624));
   INVX1 U5961 ( .A(digest[122]), .Y(n4960));
   OAI21X1 U5962 ( .A(n3082),  .B(n4962),  .C(n2425), .Y(n1623));
   INVX1 U5963 ( .A(digest[123]), .Y(n4962));
   OAI21X1 U5964 ( .A(n3083),  .B(n4964),  .C(n2360), .Y(n1622));
   AOI21X1 U5965 ( .A(N706),  .B(n3085),  .C(n3093), .Y(n4965));
   INVX1 U5966 ( .A(digest[124]), .Y(n4964));
   OAI21X1 U5967 ( .A(n4713),  .B(n4966),  .C(n2482), .Y(n1621));
   INVX1 U5968 ( .A(digest[125]), .Y(n4966));
   OAI21X1 U5969 ( .A(n3082),  .B(n4968),  .C(n2190), .Y(n1620));
   AOI21X1 U5970 ( .A(N708),  .B(n3085),  .C(n3093), .Y(n4969));
   INVX1 U5971 ( .A(digest[126]), .Y(n4968));
   OAI21X1 U5972 ( .A(n4713),  .B(n4970),  .C(n2839), .Y(n1619));
   INVX1 U5973 ( .A(digest[127]), .Y(n4970));
   OAI21X1 U5974 ( .A(n2126),  .B(n4972),  .C(n4973), .Y(n1618));
   AOI22X1 U5975 ( .A(e_reg[0]),  .B(n2977),  .C(digest[64]),  .D(n4718), .Y(n4973));
   INVX1 U5976 ( .A(f_reg[0]), .Y(n4972));
   OAI21X1 U5977 ( .A(n2126),  .B(n4974),  .C(n4975), .Y(n1617));
   AOI22X1 U5978 ( .A(e_reg[1]),  .B(n2980),  .C(digest[65]),  .D(n4718), .Y(n4975));
   INVX1 U5979 ( .A(f_reg[1]), .Y(n4974));
   NAND3X1 U5980 ( .A(n4976),  .B(n3091),  .C(n4977), .Y(n1616));
   AOI22X1 U5981 ( .A(e_reg[2]),  .B(n2978),  .C(f_reg[2]),  .D(n3088), .Y(n4977));
   NAND2X1 U5982 ( .A(digest[66]),  .B(n3038), .Y(n4976));
   NAND3X1 U5983 ( .A(n4978),  .B(n3090),  .C(n4979), .Y(n1615));
   AOI22X1 U5984 ( .A(e_reg[3]),  .B(n2977),  .C(f_reg[3]),  .D(n3088), .Y(n4979));
   NAND2X1 U5985 ( .A(digest[67]),  .B(n3027), .Y(n4978));
   OAI21X1 U5986 ( .A(n2126),  .B(n4980),  .C(n4981), .Y(n1614));
   AOI22X1 U5987 ( .A(e_reg[4]),  .B(n2978),  .C(digest[68]),  .D(n4718), .Y(n4981));
   OAI21X1 U5988 ( .A(n2126),  .B(n4982),  .C(n4983), .Y(n1613));
   AOI22X1 U5989 ( .A(e_reg[5]),  .B(n2978),  .C(digest[69]),  .D(n4718), .Y(n4983));
   INVX1 U5990 ( .A(f_reg[5]), .Y(n4982));
   OAI21X1 U5991 ( .A(n2126),  .B(n4984),  .C(n4985), .Y(n1612));
   AOI22X1 U5992 ( .A(e_reg[6]),  .B(n2977),  .C(digest[70]),  .D(n4718), .Y(n4985));
   NAND3X1 U5993 ( .A(n4986),  .B(n3091),  .C(n4987), .Y(n1611));
   AOI22X1 U5994 ( .A(e_reg[7]),  .B(n2979),  .C(f_reg[7]),  .D(n3089), .Y(n4987));
   NAND2X1 U5995 ( .A(digest[71]),  .B(n3029), .Y(n4986));
   OAI21X1 U5996 ( .A(n2126),  .B(n4988),  .C(n4989), .Y(n1610));
   AOI22X1 U5997 ( .A(e_reg[8]),  .B(n2980),  .C(digest[72]),  .D(n4718), .Y(n4989));
   INVX1 U5998 ( .A(f_reg[8]), .Y(n4988));
   OAI21X1 U5999 ( .A(n2126),  .B(n4990),  .C(n4991), .Y(n1609));
   AOI22X1 U6000 ( .A(e_reg[9]),  .B(n2980),  .C(digest[73]),  .D(n4718), .Y(n4991));
   OAI21X1 U6001 ( .A(n2126),  .B(n4992),  .C(n4993), .Y(n1608));
   AOI22X1 U6002 ( .A(e_reg[10]),  .B(n2977),  .C(digest[74]),  .D(n4718), .Y(n4993));
   NAND3X1 U6003 ( .A(n4994),  .B(n3091),  .C(n4995), .Y(n1607));
   AOI22X1 U6004 ( .A(e_reg[11]),  .B(n2979),  .C(f_reg[11]),  .D(n3089), .Y(n4995));
   NAND2X1 U6005 ( .A(digest[75]),  .B(n3036), .Y(n4994));
   OAI21X1 U6006 ( .A(n2126),  .B(n4996),  .C(n4997), .Y(n1606));
   AOI22X1 U6007 ( .A(e_reg[12]),  .B(n2977),  .C(digest[76]),  .D(n4718), .Y(n4997));
   INVX1 U6008 ( .A(f_reg[12]), .Y(n4996));
   NAND3X1 U6009 ( .A(n4998),  .B(n3090),  .C(n4999), .Y(n1605));
   AOI22X1 U6010 ( .A(e_reg[13]),  .B(n2977),  .C(f_reg[13]),  .D(n3089), .Y(n4999));
   NAND2X1 U6011 ( .A(digest[77]),  .B(n3023), .Y(n4998));
   NAND3X1 U6012 ( .A(n5000),  .B(n3090),  .C(n5001), .Y(n1604));
   AOI22X1 U6013 ( .A(e_reg[14]),  .B(n2977),  .C(f_reg[14]),  .D(n3089), .Y(n5001));
   NAND2X1 U6014 ( .A(digest[78]),  .B(n3033), .Y(n5000));
   OAI21X1 U6015 ( .A(n2126),  .B(n5002),  .C(n5003), .Y(n1603));
   AOI22X1 U6016 ( .A(e_reg[15]),  .B(n2977),  .C(digest[79]),  .D(n4718), .Y(n5003));
   INVX1 U6017 ( .A(f_reg[15]), .Y(n5002));
   NAND3X1 U6018 ( .A(n5004),  .B(n3090),  .C(n5005), .Y(n1602));
   AOI22X1 U6019 ( .A(e_reg[16]),  .B(n2977),  .C(f_reg[16]),  .D(n3088), .Y(n5005));
   NAND2X1 U6020 ( .A(digest[80]),  .B(n3017), .Y(n5004));
   OAI21X1 U6021 ( .A(n2126),  .B(n5006),  .C(n5007), .Y(n1601));
   AOI22X1 U6022 ( .A(e_reg[17]),  .B(n2977),  .C(digest[81]),  .D(n4718), .Y(n5007));
   INVX1 U6023 ( .A(f_reg[17]), .Y(n5006));
   NAND3X1 U6024 ( .A(n5008),  .B(n3090),  .C(n5009), .Y(n1600));
   AOI22X1 U6025 ( .A(e_reg[18]),  .B(n2977),  .C(f_reg[18]),  .D(n3088), .Y(n5009));
   NAND2X1 U6026 ( .A(digest[82]),  .B(n3042), .Y(n5008));
   OAI21X1 U6027 ( .A(n2126),  .B(n5010),  .C(n5011), .Y(n1599));
   AOI22X1 U6028 ( .A(e_reg[19]),  .B(n2977),  .C(digest[83]),  .D(n4718), .Y(n5011));
   OAI21X1 U6029 ( .A(n2126),  .B(n5012),  .C(n5013), .Y(n1598));
   AOI22X1 U6030 ( .A(e_reg[20]),  .B(n2977),  .C(digest[84]),  .D(n4718), .Y(n5013));
   OAI21X1 U6031 ( .A(n2126),  .B(n5014),  .C(n5015), .Y(n1597));
   AOI22X1 U6032 ( .A(e_reg[21]),  .B(n2977),  .C(digest[85]),  .D(n4718), .Y(n5015));
   OAI21X1 U6033 ( .A(n2126),  .B(n5016),  .C(n5017), .Y(n1596));
   AOI22X1 U6034 ( .A(e_reg[22]),  .B(n2977),  .C(digest[86]),  .D(n4718), .Y(n5017));
   OAI21X1 U6035 ( .A(n2126),  .B(n5018),  .C(n5019), .Y(n1595));
   AOI22X1 U6036 ( .A(e_reg[23]),  .B(n2977),  .C(digest[87]),  .D(n4718), .Y(n5019));
   INVX1 U6037 ( .A(f_reg[23]), .Y(n5018));
   NAND3X1 U6038 ( .A(n5020),  .B(n3091),  .C(n5021), .Y(n1594));
   AOI22X1 U6039 ( .A(e_reg[24]),  .B(n2977),  .C(f_reg[24]),  .D(n3089), .Y(n5021));
   NAND2X1 U6040 ( .A(digest[88]),  .B(n3031), .Y(n5020));
   NAND3X1 U6041 ( .A(n5022),  .B(n3090),  .C(n5023), .Y(n1593));
   AOI22X1 U6042 ( .A(e_reg[25]),  .B(n2977),  .C(f_reg[25]),  .D(n3088), .Y(n5023));
   NAND2X1 U6043 ( .A(digest[89]),  .B(n3047), .Y(n5022));
   OAI21X1 U6044 ( .A(n2126),  .B(n5024),  .C(n5025), .Y(n1592));
   AOI22X1 U6045 ( .A(e_reg[26]),  .B(n2980),  .C(digest[90]),  .D(n4718), .Y(n5025));
   INVX1 U6046 ( .A(f_reg[26]), .Y(n5024));
   NAND3X1 U6047 ( .A(n5026),  .B(n3091),  .C(n5027), .Y(n1591));
   AOI22X1 U6048 ( .A(e_reg[27]),  .B(n2978),  .C(f_reg[27]),  .D(n3089), .Y(n5027));
   NAND2X1 U6049 ( .A(digest[91]),  .B(n3047), .Y(n5026));
   NAND3X1 U6050 ( .A(n5028),  .B(n3090),  .C(n5029), .Y(n1590));
   AOI22X1 U6051 ( .A(e_reg[28]),  .B(n2978),  .C(f_reg[28]),  .D(n3089), .Y(n5029));
   NAND2X1 U6052 ( .A(digest[92]),  .B(n3047), .Y(n5028));
   OAI21X1 U6053 ( .A(n2126),  .B(n5030),  .C(n5031), .Y(n1589));
   AOI22X1 U6054 ( .A(e_reg[29]),  .B(n2977),  .C(digest[93]),  .D(n4718), .Y(n5031));
   OAI21X1 U6055 ( .A(n2126),  .B(n5032),  .C(n5033), .Y(n1588));
   AOI22X1 U6056 ( .A(e_reg[30]),  .B(n2979),  .C(digest[94]),  .D(n4718), .Y(n5033));
   NAND3X1 U6057 ( .A(n5034),  .B(n3091),  .C(n5035), .Y(n1587));
   AOI22X1 U6058 ( .A(e_reg[31]),  .B(n2977),  .C(f_reg[31]),  .D(n3089), .Y(n5035));
   NAND2X1 U6059 ( .A(digest[95]),  .B(n3047), .Y(n5034));
   OAI21X1 U6060 ( .A(n3083),  .B(n5036),  .C(n2539), .Y(n1586));
   INVX1 U6061 ( .A(digest[64]), .Y(n5036));
   OAI21X1 U6062 ( .A(n4713),  .B(n5038),  .C(n2596), .Y(n1585));
   INVX1 U6063 ( .A(digest[65]), .Y(n5038));
   OAI21X1 U6064 ( .A(n3082),  .B(n5040),  .C(n2216), .Y(n1584));
   AOI21X1 U6065 ( .A(N712),  .B(n3087),  .C(n3093), .Y(n5041));
   INVX1 U6066 ( .A(digest[66]), .Y(n5040));
   OAI21X1 U6067 ( .A(n3082),  .B(n5042),  .C(n2416), .Y(n1583));
   AOI21X1 U6068 ( .A(N713),  .B(n3087),  .C(n3093), .Y(n5043));
   INVX1 U6069 ( .A(digest[67]), .Y(n5042));
   OAI21X1 U6070 ( .A(n3083),  .B(n5044),  .C(n2265), .Y(n1582));
   INVX1 U6071 ( .A(digest[68]), .Y(n5044));
   OAI21X1 U6072 ( .A(n4713),  .B(n5046),  .C(n2130), .Y(n1581));
   INVX1 U6073 ( .A(digest[69]), .Y(n5046));
   OAI21X1 U6074 ( .A(n4713),  .B(n5048),  .C(n2140), .Y(n1580));
   INVX1 U6075 ( .A(digest[70]), .Y(n5048));
   OAI21X1 U6076 ( .A(n3082),  .B(n5050),  .C(n2525), .Y(n1579));
   AOI21X1 U6077 ( .A(N717),  .B(n3085),  .C(n3093), .Y(n5051));
   INVX1 U6078 ( .A(digest[71]), .Y(n5050));
   OAI21X1 U6079 ( .A(n3082),  .B(n5052),  .C(n2153), .Y(n1578));
   INVX1 U6080 ( .A(digest[72]), .Y(n5052));
   OAI21X1 U6081 ( .A(n4713),  .B(n5054),  .C(n2172), .Y(n1577));
   INVX1 U6082 ( .A(digest[73]), .Y(n5054));
   OAI21X1 U6083 ( .A(n3082),  .B(n5056),  .C(n2369), .Y(n1576));
   INVX1 U6084 ( .A(digest[74]), .Y(n5056));
   OAI21X1 U6085 ( .A(n4713),  .B(n5058),  .C(n2583), .Y(n1575));
   AOI21X1 U6086 ( .A(N721),  .B(n3085),  .C(n3093), .Y(n5059));
   INVX1 U6087 ( .A(digest[75]), .Y(n5058));
   OAI21X1 U6088 ( .A(n3083),  .B(n5060),  .C(n2315), .Y(n1574));
   INVX1 U6089 ( .A(digest[76]), .Y(n5060));
   OAI21X1 U6090 ( .A(n3082),  .B(n5062),  .C(n2640), .Y(n1573));
   AOI21X1 U6091 ( .A(N723),  .B(n3085),  .C(n3093), .Y(n5063));
   INVX1 U6092 ( .A(digest[77]), .Y(n5062));
   OAI21X1 U6093 ( .A(n4713),  .B(n5064),  .C(n2702), .Y(n1572));
   AOI21X1 U6094 ( .A(N724),  .B(n3085),  .C(n3093), .Y(n5065));
   INVX1 U6095 ( .A(digest[78]), .Y(n5064));
   OAI21X1 U6096 ( .A(n3082),  .B(n5066),  .C(n2426), .Y(n1571));
   INVX1 U6097 ( .A(digest[79]), .Y(n5066));
   OAI21X1 U6098 ( .A(n4713),  .B(n5068),  .C(n2471), .Y(n1570));
   AOI21X1 U6099 ( .A(N726),  .B(n3087),  .C(n3093), .Y(n5069));
   INVX1 U6100 ( .A(digest[80]), .Y(n5068));
   OAI21X1 U6101 ( .A(n3082),  .B(n5070),  .C(n2222), .Y(n1569));
   INVX1 U6102 ( .A(digest[81]), .Y(n5070));
   OAI21X1 U6103 ( .A(n3083),  .B(n5072),  .C(n2766), .Y(n1568));
   AOI21X1 U6104 ( .A(N728),  .B(n3085),  .C(n3093), .Y(n5073));
   INVX1 U6105 ( .A(digest[82]), .Y(n5072));
   OAI21X1 U6106 ( .A(n4713),  .B(n5074),  .C(n2540), .Y(n1567));
   INVX1 U6107 ( .A(digest[83]), .Y(n5074));
   OAI21X1 U6108 ( .A(n3082),  .B(n5076),  .C(n2658), .Y(n1566));
   INVX1 U6109 ( .A(digest[84]), .Y(n5076));
   OAI21X1 U6110 ( .A(n3083),  .B(n5078),  .C(n2131), .Y(n1565));
   INVX1 U6111 ( .A(digest[85]), .Y(n5078));
   OAI21X1 U6112 ( .A(n3082),  .B(n5080),  .C(n2141), .Y(n1564));
   INVX1 U6113 ( .A(digest[86]), .Y(n5080));
   OAI21X1 U6114 ( .A(n3083),  .B(n5082),  .C(n2154), .Y(n1563));
   INVX1 U6115 ( .A(digest[87]), .Y(n5082));
   OAI21X1 U6116 ( .A(n3082),  .B(n5084),  .C(n2829), .Y(n1562));
   AOI21X1 U6117 ( .A(N734),  .B(n3085),  .C(n3093), .Y(n5085));
   INVX1 U6118 ( .A(digest[88]), .Y(n5084));
   OAI21X1 U6119 ( .A(n3083),  .B(n5086),  .C(n2936), .Y(n1561));
   AOI21X1 U6120 ( .A(N735),  .B(n3085),  .C(n3093), .Y(n5087));
   INVX1 U6121 ( .A(digest[89]), .Y(n5086));
   OAI21X1 U6122 ( .A(n3082),  .B(n5088),  .C(n2173), .Y(n1560));
   INVX1 U6123 ( .A(digest[90]), .Y(n5088));
   OAI21X1 U6124 ( .A(n3083),  .B(n5090),  .C(n2307), .Y(n1559));
   AOI21X1 U6125 ( .A(N737),  .B(n3085),  .C(n3093), .Y(n5091));
   INVX1 U6126 ( .A(digest[91]), .Y(n5090));
   OAI21X1 U6127 ( .A(n3083),  .B(n5092),  .C(n2361), .Y(n1558));
   AOI21X1 U6128 ( .A(N738),  .B(n3085),  .C(n3093), .Y(n5093));
   INVX1 U6129 ( .A(digest[92]), .Y(n5092));
   OAI21X1 U6130 ( .A(n3083),  .B(n5094),  .C(n2194), .Y(n1557));
   INVX1 U6131 ( .A(digest[93]), .Y(n5094));
   OAI21X1 U6132 ( .A(n4713),  .B(n5096),  .C(n2223), .Y(n1556));
   INVX1 U6133 ( .A(digest[94]), .Y(n5096));
   OAI21X1 U6134 ( .A(n3082),  .B(n5098),  .C(n5099), .Y(n1555));
   AOI21X1 U6135 ( .A(N741),  .B(n3085),  .C(n4783), .Y(n5099));
   INVX1 U6136 ( .A(digest[95]), .Y(n5098));
   NAND3X1 U6137 ( .A(n5100),  .B(n3090),  .C(n5101), .Y(n1554));
   AOI22X1 U6138 ( .A(f_reg[0]),  .B(n2980),  .C(g_reg[0]),  .D(n3088), .Y(n5101));
   NAND2X1 U6139 ( .A(digest[32]),  .B(n3047), .Y(n5100));
   NAND3X1 U6140 ( .A(n5102),  .B(n3091),  .C(n5103), .Y(n1553));
   AOI22X1 U6141 ( .A(f_reg[1]),  .B(n2977),  .C(g_reg[1]),  .D(n3088), .Y(n5103));
   NAND2X1 U6142 ( .A(digest[33]),  .B(n3047), .Y(n5102));
   OAI21X1 U6143 ( .A(n2126),  .B(n5104),  .C(n5105), .Y(n1552));
   AOI22X1 U6144 ( .A(f_reg[2]),  .B(n2979),  .C(digest[34]),  .D(n4718), .Y(n5105));
   INVX1 U6145 ( .A(g_reg[2]), .Y(n5104));
   NAND3X1 U6146 ( .A(n5106),  .B(n3090),  .C(n5107), .Y(n1551));
   AOI22X1 U6147 ( .A(f_reg[3]),  .B(n2978),  .C(g_reg[3]),  .D(n3089), .Y(n5107));
   NAND2X1 U6148 ( .A(digest[35]),  .B(n3047), .Y(n5106));
   OAI21X1 U6149 ( .A(n2126),  .B(n5108),  .C(n5109), .Y(n1550));
   AOI22X1 U6150 ( .A(f_reg[4]),  .B(n2979),  .C(digest[36]),  .D(n4718), .Y(n5109));
   NAND3X1 U6151 ( .A(n5110),  .B(n3091),  .C(n5111), .Y(n1549));
   AOI22X1 U6152 ( .A(f_reg[5]),  .B(n2979),  .C(g_reg[5]),  .D(n3089), .Y(n5111));
   NAND2X1 U6153 ( .A(digest[37]),  .B(n3047), .Y(n5110));
   OAI21X1 U6154 ( .A(n2126),  .B(n5112),  .C(n5113), .Y(n1548));
   AOI22X1 U6155 ( .A(f_reg[6]),  .B(n2978),  .C(digest[38]),  .D(n4718), .Y(n5113));
   NAND3X1 U6156 ( .A(n5114),  .B(n3090),  .C(n5115), .Y(n1547));
   AOI22X1 U6157 ( .A(f_reg[7]),  .B(n2978),  .C(g_reg[7]),  .D(n3089), .Y(n5115));
   NAND2X1 U6158 ( .A(digest[39]),  .B(n3047), .Y(n5114));
   NAND3X1 U6159 ( .A(n5116),  .B(n3091),  .C(n5117), .Y(n1546));
   AOI22X1 U6160 ( .A(f_reg[8]),  .B(n2980),  .C(g_reg[8]),  .D(n3088), .Y(n5117));
   NAND2X1 U6161 ( .A(digest[40]),  .B(n3047), .Y(n5116));
   OAI21X1 U6162 ( .A(n2126),  .B(n5118),  .C(n5119), .Y(n1545));
   AOI22X1 U6163 ( .A(f_reg[9]),  .B(n2979),  .C(digest[41]),  .D(n4718), .Y(n5119));
   OAI21X1 U6164 ( .A(n2126),  .B(n5120),  .C(n5121), .Y(n1544));
   AOI22X1 U6165 ( .A(f_reg[10]),  .B(n2977),  .C(digest[42]),  .D(n4718), .Y(n5121));
   NAND3X1 U6166 ( .A(n5122),  .B(n3090),  .C(n5123), .Y(n1543));
   AOI22X1 U6167 ( .A(f_reg[11]),  .B(n2978),  .C(g_reg[11]),  .D(n3088), .Y(n5123));
   NAND2X1 U6168 ( .A(digest[43]),  .B(n3047), .Y(n5122));
   NAND3X1 U6169 ( .A(n5124),  .B(n3091),  .C(n5125), .Y(n1542));
   AOI22X1 U6170 ( .A(f_reg[12]),  .B(n2978),  .C(g_reg[12]),  .D(n3088), .Y(n5125));
   NAND2X1 U6171 ( .A(digest[44]),  .B(n3047), .Y(n5124));
   OAI21X1 U6172 ( .A(n2126),  .B(n5126),  .C(n5127), .Y(n1541));
   AOI22X1 U6173 ( .A(f_reg[13]),  .B(n2980),  .C(digest[45]),  .D(n4718), .Y(n5127));
   INVX1 U6174 ( .A(g_reg[13]), .Y(n5126));
   NAND3X1 U6175 ( .A(n5128),  .B(n3090),  .C(n5129), .Y(n1540));
   AOI22X1 U6176 ( .A(f_reg[14]),  .B(n2980),  .C(g_reg[14]),  .D(n3089), .Y(n5129));
   NAND2X1 U6177 ( .A(digest[46]),  .B(n3047), .Y(n5128));
   NAND3X1 U6178 ( .A(n5130),  .B(n3091),  .C(n5131), .Y(n1539));
   AOI22X1 U6179 ( .A(f_reg[15]),  .B(n2979),  .C(g_reg[15]),  .D(n3088), .Y(n5131));
   NAND2X1 U6180 ( .A(digest[47]),  .B(n3047), .Y(n5130));
   NAND3X1 U6181 ( .A(n5132),  .B(n3090),  .C(n5133), .Y(n1538));
   AOI22X1 U6182 ( .A(f_reg[16]),  .B(n2977),  .C(g_reg[16]),  .D(n3089), .Y(n5133));
   NAND2X1 U6183 ( .A(digest[48]),  .B(n3047), .Y(n5132));
   NAND3X1 U6184 ( .A(n5134),  .B(n3090),  .C(n5135), .Y(n1537));
   AOI22X1 U6185 ( .A(f_reg[17]),  .B(n2980),  .C(g_reg[17]),  .D(n3088), .Y(n5135));
   NAND2X1 U6186 ( .A(digest[49]),  .B(n3047), .Y(n5134));
   OAI21X1 U6187 ( .A(n2126),  .B(n5136),  .C(n5137), .Y(n1536));
   AOI22X1 U6188 ( .A(f_reg[18]),  .B(n2978),  .C(digest[50]),  .D(n4718), .Y(n5137));
   INVX1 U6189 ( .A(g_reg[18]), .Y(n5136));
   OAI21X1 U6190 ( .A(n2126),  .B(n5138),  .C(n5139), .Y(n1535));
   AOI22X1 U6191 ( .A(f_reg[19]),  .B(n2979),  .C(digest[51]),  .D(n4718), .Y(n5139));
   OAI21X1 U6192 ( .A(n2126),  .B(n5140),  .C(n5141), .Y(n1534));
   AOI22X1 U6193 ( .A(f_reg[20]),  .B(n2980),  .C(digest[52]),  .D(n4718), .Y(n5141));
   OAI21X1 U6194 ( .A(n2126),  .B(n5142),  .C(n5143), .Y(n1533));
   AOI22X1 U6195 ( .A(f_reg[21]),  .B(n2980),  .C(digest[53]),  .D(n4718), .Y(n5143));
   OAI21X1 U6196 ( .A(n2126),  .B(n5144),  .C(n5145), .Y(n1532));
   AOI22X1 U6197 ( .A(f_reg[22]),  .B(n2977),  .C(digest[54]),  .D(n4718), .Y(n5145));
   NAND3X1 U6198 ( .A(n5146),  .B(n3091),  .C(n5147), .Y(n1531));
   AOI22X1 U6199 ( .A(f_reg[23]),  .B(n2980),  .C(g_reg[23]),  .D(n3089), .Y(n5147));
   NAND2X1 U6200 ( .A(digest[55]),  .B(n3047), .Y(n5146));
   NAND3X1 U6201 ( .A(n5148),  .B(n3090),  .C(n5149), .Y(n1530));
   AOI22X1 U6202 ( .A(f_reg[24]),  .B(n2978),  .C(g_reg[24]),  .D(n3088), .Y(n5149));
   NAND2X1 U6203 ( .A(digest[56]),  .B(n3046), .Y(n5148));
   NAND3X1 U6204 ( .A(n5150),  .B(n3091),  .C(n5151), .Y(n1529));
   AOI22X1 U6205 ( .A(f_reg[25]),  .B(n2980),  .C(g_reg[25]),  .D(n3089), .Y(n5151));
   NAND2X1 U6206 ( .A(digest[57]),  .B(n3046), .Y(n5150));
   NAND3X1 U6207 ( .A(n5152),  .B(n3091),  .C(n5153), .Y(n1528));
   AOI22X1 U6208 ( .A(f_reg[26]),  .B(n2978),  .C(g_reg[26]),  .D(n3088), .Y(n5153));
   NAND2X1 U6209 ( .A(digest[58]),  .B(n3046), .Y(n5152));
   NAND3X1 U6210 ( .A(n5154),  .B(n3090),  .C(n5155), .Y(n1527));
   AOI22X1 U6211 ( .A(f_reg[27]),  .B(n2980),  .C(g_reg[27]),  .D(n3089), .Y(n5155));
   NAND2X1 U6212 ( .A(digest[59]),  .B(n3046), .Y(n5154));
   NAND3X1 U6213 ( .A(n5156),  .B(n3090),  .C(n5157), .Y(n1526));
   AOI22X1 U6214 ( .A(f_reg[28]),  .B(n2980),  .C(g_reg[28]),  .D(n3088), .Y(n5157));
   NAND2X1 U6215 ( .A(digest[60]),  .B(n3046), .Y(n5156));
   OAI21X1 U6216 ( .A(n2126),  .B(n5158),  .C(n5159), .Y(n1525));
   AOI22X1 U6217 ( .A(f_reg[29]),  .B(n2979),  .C(digest[61]),  .D(n4718), .Y(n5159));
   OAI21X1 U6218 ( .A(n2126),  .B(n5160),  .C(n5161), .Y(n1524));
   AOI22X1 U6219 ( .A(f_reg[30]),  .B(n2980),  .C(digest[62]),  .D(n4718), .Y(n5161));
   OAI21X1 U6220 ( .A(n2126),  .B(n5162),  .C(n5163), .Y(n1523));
   AOI22X1 U6221 ( .A(f_reg[31]),  .B(n2980),  .C(digest[63]),  .D(n4718), .Y(n5163));
   INVX1 U6222 ( .A(g_reg[31]), .Y(n5162));
   OAI21X1 U6223 ( .A(n4713),  .B(n5164),  .C(n5165), .Y(n1522));
   AOI21X1 U6224 ( .A(N742),  .B(n3085),  .C(n3093), .Y(n5165));
   INVX1 U6225 ( .A(digest[32]), .Y(n5164));
   OAI21X1 U6226 ( .A(n3083),  .B(n5166),  .C(n2417), .Y(n1521));
   AOI21X1 U6227 ( .A(N743),  .B(n3085),  .C(n3093), .Y(n5167));
   INVX1 U6228 ( .A(digest[33]), .Y(n5166));
   OAI21X1 U6229 ( .A(n4713),  .B(n5168),  .C(n2266), .Y(n1520));
   INVX1 U6230 ( .A(digest[34]), .Y(n5168));
   OAI21X1 U6231 ( .A(n3082),  .B(n5170),  .C(n2472), .Y(n1519));
   AOI21X1 U6232 ( .A(N745),  .B(n3085),  .C(n4783), .Y(n5171));
   INVX1 U6233 ( .A(digest[35]), .Y(n5170));
   OAI21X1 U6234 ( .A(n3082),  .B(n5172),  .C(n2597), .Y(n1518));
   INVX1 U6235 ( .A(digest[36]), .Y(n5172));
   OAI21X1 U6236 ( .A(n3083),  .B(n5174),  .C(n2526), .Y(n1517));
   AOI21X1 U6237 ( .A(N747),  .B(n3087),  .C(n3093), .Y(n5175));
   INVX1 U6238 ( .A(digest[37]), .Y(n5174));
   OAI21X1 U6239 ( .A(n4713),  .B(n5176),  .C(n2897), .Y(n1516));
   INVX1 U6240 ( .A(digest[38]), .Y(n5176));
   OAI21X1 U6241 ( .A(n3082),  .B(n5178),  .C(n2584), .Y(n1515));
   AOI21X1 U6242 ( .A(N749),  .B(n3086),  .C(n3093), .Y(n5179));
   INVX1 U6243 ( .A(digest[39]), .Y(n5178));
   OAI21X1 U6244 ( .A(n3082),  .B(n5180),  .C(n2641), .Y(n1514));
   AOI21X1 U6245 ( .A(N750),  .B(n3085),  .C(n4783), .Y(n5181));
   INVX1 U6246 ( .A(digest[40]), .Y(n5180));
   OAI21X1 U6247 ( .A(n3082),  .B(n5182),  .C(n2316), .Y(n1513));
   INVX1 U6248 ( .A(digest[41]), .Y(n5182));
   OAI21X1 U6249 ( .A(n3082),  .B(n5184),  .C(n2370), .Y(n1512));
   INVX1 U6250 ( .A(digest[42]), .Y(n5184));
   OAI21X1 U6251 ( .A(n3082),  .B(n5186),  .C(n2703), .Y(n1511));
   AOI21X1 U6252 ( .A(N753),  .B(n3086),  .C(n4783), .Y(n5187));
   INVX1 U6253 ( .A(digest[43]), .Y(n5186));
   OAI21X1 U6254 ( .A(n3082),  .B(n5188),  .C(n2767), .Y(n1510));
   AOI21X1 U6255 ( .A(N754),  .B(n3085),  .C(n3093), .Y(n5189));
   INVX1 U6256 ( .A(digest[44]), .Y(n5188));
   OAI21X1 U6257 ( .A(n3082),  .B(n5190),  .C(n2427), .Y(n1509));
   INVX1 U6258 ( .A(digest[45]), .Y(n5190));
   OAI21X1 U6259 ( .A(n3082),  .B(n5192),  .C(n2830), .Y(n1508));
   AOI21X1 U6260 ( .A(N756),  .B(n3086),  .C(n4783), .Y(n5193));
   INVX1 U6261 ( .A(digest[46]), .Y(n5192));
   OAI21X1 U6262 ( .A(n3082),  .B(n5194),  .C(n2937), .Y(n1507));
   AOI21X1 U6263 ( .A(N757),  .B(n3085),  .C(n3093), .Y(n5195));
   INVX1 U6264 ( .A(digest[47]), .Y(n5194));
   OAI21X1 U6265 ( .A(n3082),  .B(n5196),  .C(n2258), .Y(n1506));
   AOI21X1 U6266 ( .A(N758),  .B(n3087),  .C(n3093), .Y(n5197));
   INVX1 U6267 ( .A(digest[48]), .Y(n5196));
   OAI21X1 U6268 ( .A(n3082),  .B(n5198),  .C(n2308), .Y(n1505));
   AOI21X1 U6269 ( .A(N759),  .B(n3086),  .C(n3093), .Y(n5199));
   INVX1 U6270 ( .A(digest[49]), .Y(n5198));
   OAI21X1 U6271 ( .A(n3082),  .B(n5200),  .C(n2483), .Y(n1504));
   INVX1 U6272 ( .A(digest[50]), .Y(n5200));
   OAI21X1 U6273 ( .A(n3082),  .B(n5202),  .C(n2541), .Y(n1503));
   INVX1 U6274 ( .A(digest[51]), .Y(n5202));
   OAI21X1 U6275 ( .A(n4713),  .B(n5204),  .C(n2659), .Y(n1502));
   INVX1 U6276 ( .A(digest[52]), .Y(n5204));
   OAI21X1 U6277 ( .A(n4713),  .B(n5206),  .C(n2722), .Y(n1501));
   INVX1 U6278 ( .A(digest[53]), .Y(n5206));
   OAI21X1 U6279 ( .A(n4713),  .B(n5208),  .C(n2786), .Y(n1500));
   INVX1 U6280 ( .A(digest[54]), .Y(n5208));
   OAI21X1 U6281 ( .A(n4713),  .B(n5210),  .C(n2362), .Y(n1499));
   AOI21X1 U6282 ( .A(N765),  .B(n3087),  .C(n4783), .Y(n5211));
   INVX1 U6283 ( .A(digest[55]), .Y(n5210));
   OAI21X1 U6284 ( .A(n4713),  .B(n5212),  .C(n2418), .Y(n1498));
   AOI21X1 U6285 ( .A(N766),  .B(n3087),  .C(n3093), .Y(n5213));
   INVX1 U6286 ( .A(digest[56]), .Y(n5212));
   OAI21X1 U6287 ( .A(n4713),  .B(n5214),  .C(n2473), .Y(n1497));
   AOI21X1 U6288 ( .A(N767),  .B(n3087),  .C(n4783), .Y(n5215));
   INVX1 U6289 ( .A(digest[57]), .Y(n5214));
   OAI21X1 U6290 ( .A(n4713),  .B(n5216),  .C(n2527), .Y(n1496));
   AOI21X1 U6291 ( .A(N768),  .B(n3087),  .C(n4783), .Y(n5217));
   INVX1 U6292 ( .A(digest[58]), .Y(n5216));
   OAI21X1 U6293 ( .A(n3082),  .B(n5218),  .C(n2585), .Y(n1495));
   AOI21X1 U6294 ( .A(N769),  .B(n3085),  .C(n3093), .Y(n5219));
   INVX1 U6295 ( .A(digest[59]), .Y(n5218));
   OAI21X1 U6296 ( .A(n3082),  .B(n5220),  .C(n2642), .Y(n1494));
   AOI21X1 U6297 ( .A(N770),  .B(n3085),  .C(n3093), .Y(n5221));
   INVX1 U6298 ( .A(digest[60]), .Y(n5220));
   OAI21X1 U6299 ( .A(n4713),  .B(n5222),  .C(n2132), .Y(n1493));
   INVX1 U6300 ( .A(digest[61]), .Y(n5222));
   OAI21X1 U6301 ( .A(n3083),  .B(n5224),  .C(n2142), .Y(n1492));
   INVX1 U6302 ( .A(digest[62]), .Y(n5224));
   OAI21X1 U6303 ( .A(n4713),  .B(n5226),  .C(n2946), .Y(n1491));
   INVX1 U6304 ( .A(digest[63]), .Y(n5226));
   NAND3X1 U6305 ( .A(n5228),  .B(n3091),  .C(n5229), .Y(n1490));
   AOI22X1 U6306 ( .A(g_reg[0]),  .B(n2980),  .C(h_reg[0]),  .D(n3089), .Y(n5229));
   NAND2X1 U6307 ( .A(digest[0]),  .B(n3046), .Y(n5228));
   NAND2X1 U6308 ( .A(n5230),  .B(n5231), .Y(n1489));
   NAND2X1 U6309 ( .A(h_reg[1]),  .B(n3089), .Y(n5231));
   AOI22X1 U6310 ( .A(g_reg[1]),  .B(n2980),  .C(digest[1]),  .D(n4718), .Y(n5230));
   NAND2X1 U6311 ( .A(n5232),  .B(n5233), .Y(n1488));
   NAND2X1 U6312 ( .A(h_reg[2]),  .B(n3089), .Y(n5233));
   AOI22X1 U6313 ( .A(g_reg[2]),  .B(n2980),  .C(digest[2]),  .D(n4718), .Y(n5232));
   NAND3X1 U6314 ( .A(n5234),  .B(n3090),  .C(n5235), .Y(n1487));
   AOI22X1 U6315 ( .A(g_reg[3]),  .B(n2980),  .C(h_reg[3]),  .D(n3088), .Y(n5235));
   NAND2X1 U6316 ( .A(digest[3]),  .B(n3046), .Y(n5234));
   NAND3X1 U6317 ( .A(n5236),  .B(n3091),  .C(n5237), .Y(n1486));
   AOI22X1 U6318 ( .A(g_reg[4]),  .B(n2980),  .C(h_reg[4]),  .D(n3089), .Y(n5237));
   NAND2X1 U6319 ( .A(digest[4]),  .B(n3046), .Y(n5236));
   NAND2X1 U6320 ( .A(n5238),  .B(n5239), .Y(n1485));
   NAND2X1 U6321 ( .A(h_reg[5]),  .B(n3088), .Y(n5239));
   AOI22X1 U6322 ( .A(g_reg[5]),  .B(n2980),  .C(digest[5]),  .D(n4718), .Y(n5238));
   NAND2X1 U6323 ( .A(n5240),  .B(n5241), .Y(n1484));
   NAND2X1 U6324 ( .A(h_reg[6]),  .B(n3089), .Y(n5241));
   AOI22X1 U6325 ( .A(g_reg[6]),  .B(n2980),  .C(digest[6]),  .D(n4718), .Y(n5240));
   NAND2X1 U6326 ( .A(n5242),  .B(n5243), .Y(n1483));
   NAND2X1 U6327 ( .A(h_reg[7]),  .B(n3088), .Y(n5243));
   AOI22X1 U6328 ( .A(g_reg[7]),  .B(n2980),  .C(digest[7]),  .D(n4718), .Y(n5242));
   NAND3X1 U6329 ( .A(n5244),  .B(n3091),  .C(n5245), .Y(n1482));
   AOI22X1 U6330 ( .A(g_reg[8]),  .B(n2979),  .C(h_reg[8]),  .D(n3088), .Y(n5245));
   NAND2X1 U6331 ( .A(digest[8]),  .B(n3044), .Y(n5244));
   NAND2X1 U6332 ( .A(n5246),  .B(n5247), .Y(n1481));
   NAND2X1 U6333 ( .A(h_reg[9]),  .B(n3088), .Y(n5247));
   AOI22X1 U6334 ( .A(g_reg[9]),  .B(n2980),  .C(digest[9]),  .D(n4718), .Y(n5246));
   NAND3X1 U6335 ( .A(n5248),  .B(n3090),  .C(n5249), .Y(n1480));
   AOI22X1 U6336 ( .A(g_reg[10]),  .B(n2978),  .C(h_reg[10]),  .D(n3089), .Y(n5249));
   NAND2X1 U6337 ( .A(digest[10]),  .B(n3046), .Y(n5248));
   NAND3X1 U6338 ( .A(n5250),  .B(n3091),  .C(n5251), .Y(n1479));
   AOI22X1 U6339 ( .A(g_reg[11]),  .B(n2980),  .C(h_reg[11]),  .D(n3088), .Y(n5251));
   NAND2X1 U6340 ( .A(digest[11]),  .B(n3048), .Y(n5250));
   NAND2X1 U6341 ( .A(n5252),  .B(n5253), .Y(n1478));
   NAND2X1 U6342 ( .A(h_reg[12]),  .B(n3088), .Y(n5253));
   AOI22X1 U6343 ( .A(g_reg[12]),  .B(n2979),  .C(digest[12]),  .D(n4718), .Y(n5252));
   NAND2X1 U6344 ( .A(n5254),  .B(n5255), .Y(n1477));
   NAND2X1 U6345 ( .A(h_reg[13]),  .B(n3089), .Y(n5255));
   AOI22X1 U6346 ( .A(g_reg[13]),  .B(n2978),  .C(digest[13]),  .D(n4718), .Y(n5254));
   NAND3X1 U6347 ( .A(n5256),  .B(n3090),  .C(n5257), .Y(n1476));
   AOI22X1 U6348 ( .A(g_reg[14]),  .B(n2979),  .C(h_reg[14]),  .D(n3089), .Y(n5257));
   NAND2X1 U6349 ( .A(digest[14]),  .B(n3048), .Y(n5256));
   NAND3X1 U6350 ( .A(n5258),  .B(n3090),  .C(n5259), .Y(n1475));
   AOI22X1 U6351 ( .A(g_reg[15]),  .B(n2978),  .C(h_reg[15]),  .D(n3089), .Y(n5259));
   NAND2X1 U6352 ( .A(digest[15]),  .B(n3043), .Y(n5258));
   NAND2X1 U6353 ( .A(n5260),  .B(n5261), .Y(n1474));
   NAND2X1 U6354 ( .A(h_reg[16]),  .B(n3088), .Y(n5261));
   AOI22X1 U6355 ( .A(g_reg[16]),  .B(n2979),  .C(digest[16]),  .D(n4718), .Y(n5260));
   NAND2X1 U6356 ( .A(n5262),  .B(n5263), .Y(n1473));
   NAND2X1 U6357 ( .A(h_reg[17]),  .B(n3089), .Y(n5263));
   AOI22X1 U6358 ( .A(g_reg[17]),  .B(n2980),  .C(digest[17]),  .D(n4718), .Y(n5262));
   NAND2X1 U6359 ( .A(n5264),  .B(n5265), .Y(n1472));
   NAND2X1 U6360 ( .A(h_reg[18]),  .B(n3089), .Y(n5265));
   AOI22X1 U6361 ( .A(g_reg[18]),  .B(n2980),  .C(digest[18]),  .D(n4718), .Y(n5264));
   NAND2X1 U6362 ( .A(n5266),  .B(n5267), .Y(n1471));
   NAND2X1 U6363 ( .A(h_reg[19]),  .B(n3088), .Y(n5267));
   AOI22X1 U6364 ( .A(g_reg[19]),  .B(n2980),  .C(digest[19]),  .D(n4718), .Y(n5266));
   NAND2X1 U6365 ( .A(n5268),  .B(n5269), .Y(n1470));
   NAND2X1 U6366 ( .A(h_reg[20]),  .B(n3088), .Y(n5269));
   AOI22X1 U6367 ( .A(g_reg[20]),  .B(n2978),  .C(digest[20]),  .D(n4718), .Y(n5268));
   NAND3X1 U6368 ( .A(n5270),  .B(n3090),  .C(n5271), .Y(n1469));
   AOI22X1 U6369 ( .A(g_reg[21]),  .B(n2977),  .C(h_reg[21]),  .D(n3088), .Y(n5271));
   NAND2X1 U6370 ( .A(digest[21]),  .B(n3045), .Y(n5270));
   NAND3X1 U6371 ( .A(n5272),  .B(n3091),  .C(n5273), .Y(n1468));
   AOI22X1 U6372 ( .A(g_reg[22]),  .B(n2979),  .C(h_reg[22]),  .D(n3089), .Y(n5273));
   NAND2X1 U6373 ( .A(digest[22]),  .B(n3047), .Y(n5272));
   NAND3X1 U6374 ( .A(n5274),  .B(n3090),  .C(n5275), .Y(n1467));
   AOI22X1 U6375 ( .A(g_reg[23]),  .B(n2978),  .C(h_reg[23]),  .D(n3089), .Y(n5275));
   NAND2X1 U6376 ( .A(digest[23]),  .B(n3044), .Y(n5274));
   NAND3X1 U6377 ( .A(n5276),  .B(n3091),  .C(n5277), .Y(n1466));
   AOI22X1 U6378 ( .A(g_reg[24]),  .B(n2977),  .C(h_reg[24]),  .D(n3088), .Y(n5277));
   NAND2X1 U6379 ( .A(digest[24]),  .B(n3050), .Y(n5276));
   NAND3X1 U6380 ( .A(n5278),  .B(n3091),  .C(n5279), .Y(n1465));
   AOI22X1 U6381 ( .A(g_reg[25]),  .B(n2980),  .C(h_reg[25]),  .D(n3088), .Y(n5279));
   NAND2X1 U6382 ( .A(digest[25]),  .B(n3043), .Y(n5278));
   NAND2X1 U6383 ( .A(n5280),  .B(n5281), .Y(n1464));
   NAND2X1 U6384 ( .A(h_reg[26]),  .B(n3089), .Y(n5281));
   AOI22X1 U6385 ( .A(g_reg[26]),  .B(n2979),  .C(digest[26]),  .D(n4718), .Y(n5280));
   NAND3X1 U6386 ( .A(n5282),  .B(n3091),  .C(n5283), .Y(n1463));
   AOI22X1 U6387 ( .A(g_reg[27]),  .B(n2980),  .C(h_reg[27]),  .D(n3088), .Y(n5283));
   NAND2X1 U6388 ( .A(digest[27]),  .B(n3046), .Y(n5282));
   NAND3X1 U6389 ( .A(n5284),  .B(n3090),  .C(n5285), .Y(n1462));
   AOI22X1 U6390 ( .A(g_reg[28]),  .B(n2980),  .C(h_reg[28]),  .D(n3088), .Y(n5285));
   NAND2X1 U6391 ( .A(digest[28]),  .B(n3043), .Y(n5284));
   NAND2X1 U6392 ( .A(n5286),  .B(n5287), .Y(n1461));
   NAND2X1 U6393 ( .A(h_reg[29]),  .B(n3088), .Y(n5287));
   AOI22X1 U6394 ( .A(g_reg[29]),  .B(n2979),  .C(digest[29]),  .D(n4718), .Y(n5286));
   NAND3X1 U6395 ( .A(n5288),  .B(n3090),  .C(n5289), .Y(n1460));
   AOI22X1 U6396 ( .A(g_reg[30]),  .B(n2979),  .C(h_reg[30]),  .D(n3088), .Y(n5289));
   NAND2X1 U6397 ( .A(digest[30]),  .B(n3043), .Y(n5288));
   NAND2X1 U6398 ( .A(n5290),  .B(n5291), .Y(n1459));
   NAND2X1 U6399 ( .A(h_reg[31]),  .B(n3088), .Y(n5291));
   AOI22X1 U6400 ( .A(g_reg[31]),  .B(n2978),  .C(digest[31]),  .D(n4718), .Y(n5290));
   OAI21X1 U6401 ( .A(n4713),  .B(n5292),  .C(n5293), .Y(n1458));
   AOI21X1 U6402 ( .A(N774),  .B(n3087),  .C(n4783), .Y(n5293));
   INVX1 U6403 ( .A(digest[0]), .Y(n5292));
   OAI21X1 U6404 ( .A(n4713),  .B(n5294),  .C(n2155), .Y(n1457));
   INVX1 U6405 ( .A(digest[1]), .Y(n5294));
   OAI21X1 U6406 ( .A(n4713),  .B(n5296),  .C(n2174), .Y(n1456));
   INVX1 U6407 ( .A(digest[2]), .Y(n5296));
   OAI21X1 U6408 ( .A(n4713),  .B(n5298),  .C(n2704), .Y(n1455));
   AOI21X1 U6409 ( .A(N777),  .B(n3086),  .C(n3093), .Y(n5299));
   INVX1 U6410 ( .A(digest[3]), .Y(n5298));
   OAI21X1 U6411 ( .A(n3083),  .B(n5300),  .C(n2768), .Y(n1454));
   AOI21X1 U6412 ( .A(N778),  .B(n3085),  .C(n4783), .Y(n5301));
   INVX1 U6413 ( .A(digest[4]), .Y(n5300));
   OAI21X1 U6414 ( .A(n4713),  .B(n5302),  .C(n2195), .Y(n1453));
   INVX1 U6415 ( .A(digest[5]), .Y(n5302));
   OAI21X1 U6416 ( .A(n3082),  .B(n5304),  .C(n2371), .Y(n1452));
   INVX1 U6417 ( .A(digest[6]), .Y(n5304));
   OAI21X1 U6418 ( .A(n3083),  .B(n5306),  .C(n2428), .Y(n1451));
   INVX1 U6419 ( .A(digest[7]), .Y(n5306));
   OAI21X1 U6420 ( .A(n3083),  .B(n5308),  .C(n2831), .Y(n1450));
   AOI21X1 U6421 ( .A(N782),  .B(n3087),  .C(n4783), .Y(n5309));
   INVX1 U6422 ( .A(digest[8]), .Y(n5308));
   OAI21X1 U6423 ( .A(n4713),  .B(n5310),  .C(n2484), .Y(n1449));
   INVX1 U6424 ( .A(digest[9]), .Y(n5310));
   OAI21X1 U6425 ( .A(n4713),  .B(n5312),  .C(n2938), .Y(n1448));
   AOI21X1 U6426 ( .A(N784),  .B(n3087),  .C(n3093), .Y(n5313));
   INVX1 U6427 ( .A(digest[10]), .Y(n5312));
   OAI21X1 U6428 ( .A(n3082),  .B(n5314),  .C(n2259), .Y(n1447));
   AOI21X1 U6429 ( .A(N785),  .B(n3085),  .C(n4783), .Y(n5315));
   INVX1 U6430 ( .A(digest[11]), .Y(n5314));
   OAI21X1 U6431 ( .A(n3082),  .B(n5316),  .C(n2542), .Y(n1446));
   INVX1 U6432 ( .A(digest[12]), .Y(n5316));
   OAI21X1 U6433 ( .A(n4713),  .B(n5318),  .C(n2660), .Y(n1445));
   INVX1 U6434 ( .A(digest[13]), .Y(n5318));
   OAI21X1 U6435 ( .A(n4713),  .B(n5320),  .C(n2309), .Y(n1444));
   AOI21X1 U6436 ( .A(N788),  .B(n3086),  .C(n3093), .Y(n5321));
   INVX1 U6437 ( .A(digest[14]), .Y(n5320));
   OAI21X1 U6438 ( .A(n3083),  .B(n5322),  .C(n2363), .Y(n1443));
   AOI21X1 U6439 ( .A(N789),  .B(n3086),  .C(n3093), .Y(n5323));
   INVX1 U6440 ( .A(digest[15]), .Y(n5322));
   OAI21X1 U6441 ( .A(n3082),  .B(n5324),  .C(n2224), .Y(n1442));
   INVX1 U6442 ( .A(digest[16]), .Y(n5324));
   OAI21X1 U6443 ( .A(n3083),  .B(n5326),  .C(n2267), .Y(n1441));
   INVX1 U6444 ( .A(digest[17]), .Y(n5326));
   OAI21X1 U6445 ( .A(n4713),  .B(n5328),  .C(n2317), .Y(n1440));
   INVX1 U6446 ( .A(digest[18]), .Y(n5328));
   OAI21X1 U6447 ( .A(n4713),  .B(n5330),  .C(n2598), .Y(n1439));
   INVX1 U6448 ( .A(digest[19]), .Y(n5330));
   OAI21X1 U6449 ( .A(n4713),  .B(n5332),  .C(n2723), .Y(n1438));
   INVX1 U6450 ( .A(digest[20]), .Y(n5332));
   OAI21X1 U6451 ( .A(n3082),  .B(n5334),  .C(n2419), .Y(n1437));
   AOI21X1 U6452 ( .A(N795),  .B(n3087),  .C(n3093), .Y(n5335));
   INVX1 U6453 ( .A(digest[21]), .Y(n5334));
   OAI21X1 U6454 ( .A(n3083),  .B(n5336),  .C(n2474), .Y(n1436));
   AOI21X1 U6455 ( .A(N796),  .B(n3086),  .C(n4783), .Y(n5337));
   INVX1 U6456 ( .A(digest[22]), .Y(n5336));
   OAI21X1 U6457 ( .A(n3083),  .B(n5338),  .C(n2528), .Y(n1435));
   AOI21X1 U6458 ( .A(N797),  .B(n3085),  .C(n3093), .Y(n5339));
   INVX1 U6459 ( .A(digest[23]), .Y(n5338));
   OAI21X1 U6460 ( .A(n4713),  .B(n5340),  .C(n2586), .Y(n1434));
   AOI21X1 U6461 ( .A(N798),  .B(n3087),  .C(n3093), .Y(n5341));
   INVX1 U6462 ( .A(digest[24]), .Y(n5340));
   OAI21X1 U6463 ( .A(n3083),  .B(n5342),  .C(n2705), .Y(n1433));
   AOI21X1 U6464 ( .A(N799),  .B(n3086),  .C(n4783), .Y(n5343));
   INVX1 U6465 ( .A(digest[25]), .Y(n5342));
   OAI21X1 U6466 ( .A(n3082),  .B(n5344),  .C(n2787), .Y(n1432));
   INVX1 U6467 ( .A(digest[26]), .Y(n5344));
   OAI21X1 U6468 ( .A(n3083),  .B(n5346),  .C(n2939), .Y(n1431));
   AOI21X1 U6469 ( .A(N801),  .B(n3087),  .C(n4783), .Y(n5347));
   INVX1 U6470 ( .A(digest[27]), .Y(n5346));
   OAI21X1 U6471 ( .A(n3082),  .B(n5348),  .C(n2643), .Y(n1430));
   AOI21X1 U6472 ( .A(N802),  .B(n3086),  .C(n4783), .Y(n5349));
   INVX1 U6473 ( .A(digest[28]), .Y(n5348));
   OAI21X1 U6474 ( .A(n3083),  .B(n5350),  .C(n5351), .Y(n1429));
   NAND2X1 U6475 ( .A(N803),  .B(n3087), .Y(n5351));
   INVX1 U6476 ( .A(digest[29]), .Y(n5350));
   OAI21X1 U6477 ( .A(n3083),  .B(n5352),  .C(n2769), .Y(n1428));
   AOI21X1 U6478 ( .A(N804),  .B(n3086),  .C(n3093), .Y(n5353));
   INVX1 U6479 ( .A(digest[30]), .Y(n5352));
   OAI21X1 U6480 ( .A(n4713),  .B(n5354),  .C(n2947), .Y(n1427));
   INVX1 U6481 ( .A(digest[31]), .Y(n5354));
   NAND3X1 U6482 ( .A(n5356),  .B(n3090),  .C(n5357), .Y(n1426));
   AOI22X1 U6483 ( .A(N1547),  .B(n2980),  .C(a_reg[0]),  .D(n3088), .Y(n5357));
   NAND2X1 U6484 ( .A(digest[224]),  .B(n3043), .Y(n5356));
   NAND3X1 U6485 ( .A(n5358),  .B(n3091),  .C(n5359), .Y(n1425));
   AOI22X1 U6486 ( .A(N1548),  .B(n2977),  .C(a_reg[1]),  .D(n3088), .Y(n5359));
   NAND2X1 U6487 ( .A(digest[225]),  .B(n3043), .Y(n5358));
   NAND3X1 U6488 ( .A(n5360),  .B(n3090),  .C(n5361), .Y(n1424));
   AOI22X1 U6489 ( .A(N1549),  .B(n2977),  .C(n3088),  .D(a_reg[2]), .Y(n5361));
   NAND2X1 U6490 ( .A(digest[226]),  .B(n3043), .Y(n5360));
   OAI21X1 U6491 ( .A(n2126),  .B(n5362),  .C(n5363), .Y(n1423));
   AOI22X1 U6492 ( .A(N1550),  .B(n2979),  .C(digest[227]),  .D(n4718), .Y(n5363));
   OAI21X1 U6493 ( .A(n2126),  .B(n5364),  .C(n5365), .Y(n1422));
   AOI22X1 U6494 ( .A(N1551),  .B(n2980),  .C(digest[228]),  .D(n4718), .Y(n5365));
   NAND3X1 U6495 ( .A(n5366),  .B(n3090),  .C(n5367), .Y(n1421));
   AOI22X1 U6496 ( .A(N1552),  .B(n2978),  .C(a_reg[5]),  .D(n3088), .Y(n5367));
   NAND2X1 U6497 ( .A(digest[229]),  .B(n3043), .Y(n5366));
   NAND3X1 U6498 ( .A(n5368),  .B(n3091),  .C(n5369), .Y(n1420));
   AOI22X1 U6499 ( .A(N1553),  .B(n2977),  .C(a_reg[6]),  .D(n3088), .Y(n5369));
   NAND2X1 U6500 ( .A(digest[230]),  .B(n3043), .Y(n5368));
   OAI21X1 U6501 ( .A(n2126),  .B(n5370),  .C(n5371), .Y(n1419));
   AOI22X1 U6502 ( .A(N1554),  .B(n2979),  .C(digest[231]),  .D(n4718), .Y(n5371));
   OAI21X1 U6503 ( .A(n2126),  .B(n5372),  .C(n5373), .Y(n1418));
   AOI22X1 U6504 ( .A(N1555),  .B(n2980),  .C(digest[232]),  .D(n4718), .Y(n5373));
   NAND3X1 U6505 ( .A(n5374),  .B(n3090),  .C(n5375), .Y(n1417));
   AOI22X1 U6506 ( .A(N1556),  .B(n2978),  .C(n3088),  .D(a_reg[9]), .Y(n5375));
   NAND2X1 U6507 ( .A(digest[233]),  .B(n3043), .Y(n5374));
   NAND3X1 U6508 ( .A(n5376),  .B(n3091),  .C(n5377), .Y(n1416));
   AOI22X1 U6509 ( .A(N1557),  .B(n2977),  .C(n3088),  .D(a_reg[10]), .Y(n5377));
   NAND2X1 U6510 ( .A(digest[234]),  .B(n3043), .Y(n5376));
   OAI21X1 U6511 ( .A(n2126),  .B(n5378),  .C(n5379), .Y(n1415));
   AOI22X1 U6512 ( .A(N1558),  .B(n2979),  .C(digest[235]),  .D(n4718), .Y(n5379));
   OAI21X1 U6513 ( .A(n2126),  .B(n5380),  .C(n5381), .Y(n1414));
   AOI22X1 U6514 ( .A(N1559),  .B(n2980),  .C(digest[236]),  .D(n4718), .Y(n5381));
   NAND3X1 U6515 ( .A(n5382),  .B(n3090),  .C(n5383), .Y(n1413));
   AOI22X1 U6516 ( .A(N1560),  .B(n2978),  .C(a_reg[13]),  .D(n3088), .Y(n5383));
   NAND2X1 U6517 ( .A(digest[237]),  .B(n3043), .Y(n5382));
   NAND3X1 U6518 ( .A(n5384),  .B(n3091),  .C(n5385), .Y(n1412));
   AOI22X1 U6519 ( .A(N1561),  .B(n2977),  .C(a_reg[14]),  .D(n3088), .Y(n5385));
   NAND2X1 U6520 ( .A(digest[238]),  .B(n3043), .Y(n5384));
   NAND3X1 U6521 ( .A(n5386),  .B(n3090),  .C(n5387), .Y(n1411));
   AOI22X1 U6522 ( .A(N1562),  .B(n2979),  .C(a_reg[15]),  .D(n3089), .Y(n5387));
   NAND2X1 U6523 ( .A(digest[239]),  .B(n3043), .Y(n5386));
   NAND3X1 U6524 ( .A(n5388),  .B(n3091),  .C(n5389), .Y(n1410));
   AOI22X1 U6525 ( .A(N1563),  .B(n2978),  .C(a_reg[16]),  .D(n3089), .Y(n5389));
   NAND2X1 U6526 ( .A(digest[240]),  .B(n3043), .Y(n5388));
   OAI21X1 U6527 ( .A(n2126),  .B(n5390),  .C(n5391), .Y(n1409));
   AOI22X1 U6528 ( .A(N1564),  .B(n2977),  .C(digest[241]),  .D(n4718), .Y(n5391));
   OAI21X1 U6529 ( .A(n2126),  .B(n5392),  .C(n5393), .Y(n1408));
   AOI22X1 U6530 ( .A(N1565),  .B(n2977),  .C(digest[242]),  .D(n4718), .Y(n5393));
   NAND3X1 U6531 ( .A(n5394),  .B(n3090),  .C(n5395), .Y(n1407));
   AOI22X1 U6532 ( .A(N1566),  .B(n2980),  .C(a_reg[19]),  .D(n3089), .Y(n5395));
   NAND2X1 U6533 ( .A(digest[243]),  .B(n3043), .Y(n5394));
   OAI21X1 U6534 ( .A(n2126),  .B(n5396),  .C(n5397), .Y(n1406));
   AOI22X1 U6535 ( .A(N1567),  .B(n2979),  .C(digest[244]),  .D(n4718), .Y(n5397));
   OAI21X1 U6536 ( .A(n2126),  .B(n5398),  .C(n5399), .Y(n1405));
   AOI22X1 U6537 ( .A(N1568),  .B(n2978),  .C(digest[245]),  .D(n4718), .Y(n5399));
   OAI21X1 U6538 ( .A(n2126),  .B(n5400),  .C(n5401), .Y(n1404));
   AOI22X1 U6539 ( .A(N1569),  .B(n2980),  .C(digest[246]),  .D(n4718), .Y(n5401));
   OAI21X1 U6540 ( .A(n2126),  .B(n5402),  .C(n5403), .Y(n1403));
   AOI22X1 U6541 ( .A(N1570),  .B(n2977),  .C(digest[247]),  .D(n4718), .Y(n5403));
   OAI21X1 U6542 ( .A(n2126),  .B(n5404),  .C(n5405), .Y(n1402));
   AOI22X1 U6543 ( .A(N1571),  .B(n2978),  .C(digest[248]),  .D(n4718), .Y(n5405));
   NAND3X1 U6544 ( .A(n5406),  .B(n3091),  .C(n5407), .Y(n1401));
   AOI22X1 U6545 ( .A(N1572),  .B(n2978),  .C(n3088),  .D(a_reg[25]), .Y(n5407));
   NAND2X1 U6546 ( .A(digest[249]),  .B(n3043), .Y(n5406));
   OAI21X1 U6547 ( .A(n2126),  .B(n5408),  .C(n5409), .Y(n1400));
   AOI22X1 U6548 ( .A(N1573),  .B(n2980),  .C(digest[250]),  .D(n4718), .Y(n5409));
   NAND3X1 U6549 ( .A(n5410),  .B(n3091),  .C(n5411), .Y(n1399));
   AOI22X1 U6550 ( .A(N1574),  .B(n2979),  .C(n3089),  .D(a_reg[27]), .Y(n5411));
   NAND2X1 U6551 ( .A(digest[251]),  .B(n3043), .Y(n5410));
   OAI21X1 U6552 ( .A(n2126),  .B(n5412),  .C(n5413), .Y(n1398));
   AOI22X1 U6553 ( .A(N1575),  .B(n2980),  .C(digest[252]),  .D(n4718), .Y(n5413));
   NAND3X1 U6554 ( .A(n5414),  .B(n3090),  .C(n5415), .Y(n1397));
   AOI22X1 U6555 ( .A(N1576),  .B(n2977),  .C(n3089),  .D(a_reg[29]), .Y(n5415));
   NAND2X1 U6556 ( .A(digest[253]),  .B(n3044), .Y(n5414));
   NAND3X1 U6557 ( .A(n5416),  .B(n3091),  .C(n5417), .Y(n1396));
   AOI22X1 U6558 ( .A(N1577),  .B(n2980),  .C(a_reg[30]),  .D(n3088), .Y(n5417));
   NAND2X1 U6559 ( .A(digest[254]),  .B(n3044), .Y(n5416));
   OAI21X1 U6560 ( .A(n2126),  .B(n5418),  .C(n5419), .Y(n1395));
   AOI22X1 U6561 ( .A(N1578),  .B(n2978),  .C(digest[255]),  .D(n4718), .Y(n5419));
   OAI21X1 U6562 ( .A(n3083),  .B(n5420),  .C(n5421), .Y(n1394));
   AOI21X1 U6563 ( .A(N550),  .B(n3086),  .C(n3093), .Y(n5421));
   INVX1 U6564 ( .A(digest[224]), .Y(n5420));
   OAI21X1 U6565 ( .A(n3083),  .B(n5422),  .C(n2832), .Y(n1393));
   AOI21X1 U6566 ( .A(N551),  .B(n3085),  .C(n4783), .Y(n5423));
   INVX1 U6567 ( .A(digest[225]), .Y(n5422));
   OAI21X1 U6568 ( .A(n4713),  .B(n5424),  .C(n2217), .Y(n1392));
   AOI21X1 U6569 ( .A(N552),  .B(n3085),  .C(n3093), .Y(n5425));
   INVX1 U6570 ( .A(digest[226]), .Y(n5424));
   OAI21X1 U6571 ( .A(n3082),  .B(n5426),  .C(n2133), .Y(n1391));
   INVX1 U6572 ( .A(digest[227]), .Y(n5426));
   OAI21X1 U6573 ( .A(n4713),  .B(n5428),  .C(n2143), .Y(n1390));
   INVX1 U6574 ( .A(digest[228]), .Y(n5428));
   OAI21X1 U6575 ( .A(n4713),  .B(n5430),  .C(n2260), .Y(n1389));
   AOI21X1 U6576 ( .A(N555),  .B(n3086),  .C(n3093), .Y(n5431));
   INVX1 U6577 ( .A(digest[229]), .Y(n5430));
   OAI21X1 U6578 ( .A(n3082),  .B(n5432),  .C(n2475), .Y(n1388));
   AOI21X1 U6579 ( .A(N556),  .B(n3087),  .C(n4783), .Y(n5433));
   INVX1 U6580 ( .A(digest[230]), .Y(n5432));
   OAI21X1 U6581 ( .A(n3083),  .B(n5434),  .C(n2156), .Y(n1387));
   INVX1 U6582 ( .A(digest[231]), .Y(n5434));
   OAI21X1 U6583 ( .A(n4713),  .B(n5436),  .C(n2175), .Y(n1386));
   INVX1 U6584 ( .A(digest[232]), .Y(n5436));
   OAI21X1 U6585 ( .A(n3083),  .B(n5438),  .C(n2706), .Y(n1385));
   AOI21X1 U6586 ( .A(N559),  .B(n3086),  .C(n3093), .Y(n5439));
   INVX1 U6587 ( .A(digest[233]), .Y(n5438));
   OAI21X1 U6588 ( .A(n4713),  .B(n5440),  .C(n2940), .Y(n1384));
   AOI21X1 U6589 ( .A(N560),  .B(n3087),  .C(n3093), .Y(n5441));
   INVX1 U6590 ( .A(digest[234]), .Y(n5440));
   OAI21X1 U6591 ( .A(n3082),  .B(n5442),  .C(n2196), .Y(n1383));
   INVX1 U6592 ( .A(digest[235]), .Y(n5442));
   OAI21X1 U6593 ( .A(n3083),  .B(n5444),  .C(n2268), .Y(n1382));
   INVX1 U6594 ( .A(digest[236]), .Y(n5444));
   OAI21X1 U6595 ( .A(n3083),  .B(n5446),  .C(n2529), .Y(n1381));
   AOI21X1 U6596 ( .A(N563),  .B(n3086),  .C(n3093), .Y(n5447));
   INVX1 U6597 ( .A(digest[237]), .Y(n5446));
   OAI21X1 U6598 ( .A(n3083),  .B(n5448),  .C(n2587), .Y(n1380));
   AOI21X1 U6599 ( .A(N564),  .B(n3085),  .C(n3093), .Y(n5449));
   INVX1 U6600 ( .A(digest[238]), .Y(n5448));
   OAI21X1 U6601 ( .A(n4713),  .B(n5450),  .C(n2644), .Y(n1379));
   AOI21X1 U6602 ( .A(N565),  .B(n3086),  .C(n4783), .Y(n5451));
   INVX1 U6603 ( .A(digest[239]), .Y(n5450));
   OAI21X1 U6604 ( .A(n3082),  .B(n5452),  .C(n2770), .Y(n1378));
   AOI21X1 U6605 ( .A(N566),  .B(n3086),  .C(n4783), .Y(n5453));
   INVX1 U6606 ( .A(digest[240]), .Y(n5452));
   OAI21X1 U6607 ( .A(n4713),  .B(n5454),  .C(n2318), .Y(n1377));
   INVX1 U6608 ( .A(digest[241]), .Y(n5454));
   OAI21X1 U6609 ( .A(n3082),  .B(n5456),  .C(n2372), .Y(n1376));
   INVX1 U6610 ( .A(digest[242]), .Y(n5456));
   OAI21X1 U6611 ( .A(n3083),  .B(n5458),  .C(n2833), .Y(n1375));
   AOI21X1 U6612 ( .A(N569),  .B(n3085),  .C(n4783), .Y(n5459));
   INVX1 U6613 ( .A(digest[243]), .Y(n5458));
   OAI21X1 U6614 ( .A(n4713),  .B(n5460),  .C(n2225), .Y(n1374));
   INVX1 U6615 ( .A(digest[244]), .Y(n5460));
   OAI21X1 U6616 ( .A(n3082),  .B(n5462),  .C(n2429), .Y(n1373));
   INVX1 U6617 ( .A(digest[245]), .Y(n5462));
   OAI21X1 U6618 ( .A(n3083),  .B(n5464),  .C(n2485), .Y(n1372));
   INVX1 U6619 ( .A(digest[246]), .Y(n5464));
   OAI21X1 U6620 ( .A(n4713),  .B(n5466),  .C(n2543), .Y(n1371));
   INVX1 U6621 ( .A(digest[247]), .Y(n5466));
   OAI21X1 U6622 ( .A(n3083),  .B(n5468),  .C(n2599), .Y(n1370));
   INVX1 U6623 ( .A(digest[248]), .Y(n5468));
   OAI21X1 U6624 ( .A(n3082),  .B(n5470),  .C(n2310), .Y(n1369));
   AOI21X1 U6625 ( .A(N575),  .B(n3086),  .C(n3093), .Y(n5471));
   INVX1 U6626 ( .A(digest[249]), .Y(n5470));
   OAI21X1 U6627 ( .A(n3083),  .B(n5472),  .C(n2661), .Y(n1368));
   INVX1 U6628 ( .A(digest[250]), .Y(n5472));
   OAI21X1 U6629 ( .A(n3083),  .B(n5474),  .C(n2364), .Y(n1367));
   AOI21X1 U6630 ( .A(N577),  .B(n3087),  .C(n3093), .Y(n5475));
   INVX1 U6631 ( .A(digest[251]), .Y(n5474));
   OAI21X1 U6632 ( .A(n4713),  .B(n5476),  .C(n2724), .Y(n1366));
   INVX1 U6633 ( .A(digest[252]), .Y(n5476));
   OAI21X1 U6634 ( .A(n4713),  .B(n5478),  .C(n2420), .Y(n1365));
   AOI21X1 U6635 ( .A(N579),  .B(n3087),  .C(n3093), .Y(n5479));
   INVX1 U6636 ( .A(digest[253]), .Y(n5478));
   OAI21X1 U6637 ( .A(n3082),  .B(n5480),  .C(n2169), .Y(n1364));
   AOI21X1 U6638 ( .A(N580),  .B(n3085),  .C(n3093), .Y(n5481));
   INVX1 U6639 ( .A(digest[254]), .Y(n5480));
   OAI21X1 U6640 ( .A(n3082),  .B(n5482),  .C(n2948), .Y(n1363));
   INVX1 U6641 ( .A(digest[255]), .Y(n5482));
   NAND3X1 U6642 ( .A(n5484),  .B(n3091),  .C(n5485), .Y(n1362));
   AOI22X1 U6643 ( .A(a_reg[0]),  .B(n2979),  .C(b_reg[0]),  .D(n3088), .Y(n5485));
   NAND2X1 U6644 ( .A(digest[192]),  .B(n3044), .Y(n5484));
   OAI21X1 U6645 ( .A(n2126),  .B(n5486),  .C(n5487), .Y(n1361));
   AOI22X1 U6646 ( .A(a_reg[1]),  .B(n2977),  .C(digest[193]),  .D(n4718), .Y(n5487));
   NAND3X1 U6647 ( .A(n5488),  .B(n3091),  .C(n5489), .Y(n1360));
   AOI22X1 U6648 ( .A(a_reg[2]),  .B(n2978),  .C(n3088),  .D(b_reg[2]), .Y(n5489));
   NAND2X1 U6649 ( .A(digest[194]),  .B(n3044), .Y(n5488));
   OAI21X1 U6650 ( .A(n2126),  .B(n5490),  .C(n5491), .Y(n1359));
   AOI22X1 U6651 ( .A(a_reg[3]),  .B(n2979),  .C(digest[195]),  .D(n4718), .Y(n5491));
   OAI21X1 U6652 ( .A(n2126),  .B(n5492),  .C(n5493), .Y(n1358));
   AOI22X1 U6653 ( .A(a_reg[4]),  .B(n2978),  .C(digest[196]),  .D(n4718), .Y(n5493));
   OAI21X1 U6654 ( .A(n2126),  .B(n5494),  .C(n5495), .Y(n1357));
   AOI22X1 U6655 ( .A(a_reg[5]),  .B(n2978),  .C(digest[197]),  .D(n4718), .Y(n5495));
   OAI21X1 U6656 ( .A(n2126),  .B(n5496),  .C(n5497), .Y(puf_12_wire_3));
   AOI22X1 U6657 ( .A(a_reg[6]),  .B(n2979),  .C(digest[198]),  .D(n4718), .Y(n5497));
   NAND3X1 U6658 ( .A(n5498),  .B(n3090),  .C(n5499), .Y(n1355));
   AOI22X1 U6659 ( .A(a_reg[7]),  .B(n2977),  .C(b_reg[7]),  .D(n3088), .Y(n5499));
   NAND2X1 U6660 ( .A(digest[199]),  .B(n3044), .Y(n5498));
   OAI21X1 U6661 ( .A(n2126),  .B(n5500),  .C(n5501), .Y(n1354));
   AOI22X1 U6662 ( .A(a_reg[8]),  .B(n2978),  .C(digest[200]),  .D(n4718), .Y(n5501));
   NAND3X1 U6663 ( .A(n5502),  .B(n3091),  .C(n5503), .Y(n1353));
   AOI22X1 U6664 ( .A(a_reg[9]),  .B(n2979),  .C(n3089),  .D(b_reg[9]), .Y(n5503));
   NAND2X1 U6665 ( .A(digest[201]),  .B(n3044), .Y(n5502));
   NAND3X1 U6666 ( .A(n5504),  .B(n3090),  .C(n5505), .Y(n1352));
   AOI22X1 U6667 ( .A(a_reg[10]),  .B(n2978),  .C(n3089),  .D(b_reg[10]), .Y(n5505));
   NAND2X1 U6668 ( .A(digest[202]),  .B(n3044), .Y(n5504));
   NAND3X1 U6669 ( .A(n5506),  .B(n3090),  .C(n5507), .Y(n1351));
   AOI22X1 U6670 ( .A(a_reg[11]),  .B(n2980),  .C(b_reg[11]),  .D(n3089), .Y(n5507));
   NAND2X1 U6671 ( .A(digest[203]),  .B(n3044), .Y(n5506));
   OAI21X1 U6672 ( .A(n2126),  .B(n5508),  .C(n5509), .Y(n1350));
   AOI22X1 U6673 ( .A(a_reg[12]),  .B(n2977),  .C(digest[204]),  .D(n4718), .Y(n5509));
   NAND3X1 U6674 ( .A(n5510),  .B(n3091),  .C(n5511), .Y(n1349));
   AOI22X1 U6675 ( .A(a_reg[13]),  .B(n2978),  .C(b_reg[13]),  .D(n3088), .Y(n5511));
   NAND2X1 U6676 ( .A(digest[205]),  .B(n3044), .Y(n5510));
   OAI21X1 U6677 ( .A(n2126),  .B(n5512),  .C(n5513), .Y(n1348));
   AOI22X1 U6678 ( .A(a_reg[14]),  .B(n2980),  .C(digest[206]),  .D(n4718), .Y(n5513));
   NAND3X1 U6679 ( .A(n5514),  .B(n3091),  .C(n5515), .Y(n1347));
   AOI22X1 U6680 ( .A(a_reg[15]),  .B(n2978),  .C(b_reg[15]),  .D(n3088), .Y(n5515));
   NAND2X1 U6681 ( .A(digest[207]),  .B(n3044), .Y(n5514));
   NAND3X1 U6682 ( .A(n5516),  .B(n3091),  .C(n5517), .Y(n1346));
   AOI22X1 U6683 ( .A(a_reg[16]),  .B(n2977),  .C(b_reg[16]),  .D(n3089), .Y(n5517));
   NAND2X1 U6684 ( .A(digest[208]),  .B(n3044), .Y(n5516));
   NAND3X1 U6685 ( .A(n5518),  .B(n3090),  .C(n5519), .Y(n1345));
   AOI22X1 U6686 ( .A(a_reg[17]),  .B(n2979),  .C(b_reg[17]),  .D(n3088), .Y(n5519));
   NAND2X1 U6687 ( .A(digest[209]),  .B(n3044), .Y(n5518));
   NAND3X1 U6688 ( .A(n5520),  .B(n3090),  .C(n5521), .Y(n1344));
   AOI22X1 U6689 ( .A(a_reg[18]),  .B(n2979),  .C(b_reg[18]),  .D(n3088), .Y(n5521));
   NAND2X1 U6690 ( .A(digest[210]),  .B(n3044), .Y(n5520));
   OAI21X1 U6691 ( .A(n2126),  .B(n5522),  .C(n5523), .Y(n1343));
   AOI22X1 U6692 ( .A(a_reg[19]),  .B(n2978),  .C(digest[211]),  .D(n4718), .Y(n5523));
   OAI21X1 U6693 ( .A(n2126),  .B(n5524),  .C(n5525), .Y(n1342));
   AOI22X1 U6694 ( .A(a_reg[20]),  .B(n2980),  .C(digest[212]),  .D(n4718), .Y(n5525));
   NAND3X1 U6695 ( .A(n5526),  .B(n3090),  .C(n5527), .Y(n1341));
   AOI22X1 U6696 ( .A(a_reg[21]),  .B(n2977),  .C(b_reg[21]),  .D(n3088), .Y(n5527));
   NAND2X1 U6697 ( .A(digest[213]),  .B(n3044), .Y(n5526));
   NAND3X1 U6698 ( .A(n5528),  .B(n3091),  .C(n5529), .Y(n1340));
   AOI22X1 U6699 ( .A(a_reg[22]),  .B(n2977),  .C(b_reg[22]),  .D(n3088), .Y(n5529));
   NAND2X1 U6700 ( .A(digest[214]),  .B(n3044), .Y(n5528));
   OAI21X1 U6701 ( .A(n2126),  .B(n5530),  .C(n5531), .Y(n1339));
   AOI22X1 U6702 ( .A(a_reg[23]),  .B(n2977),  .C(digest[215]),  .D(n4718), .Y(n5531));
   NAND3X1 U6703 ( .A(n5532),  .B(n3091),  .C(n5533), .Y(n1338));
   AOI22X1 U6704 ( .A(a_reg[24]),  .B(n2980),  .C(b_reg[24]),  .D(n3088), .Y(n5533));
   NAND2X1 U6705 ( .A(digest[216]),  .B(n3044), .Y(n5532));
   NAND3X1 U6706 ( .A(n5534),  .B(n3091),  .C(n5535), .Y(n1337));
   AOI22X1 U6707 ( .A(a_reg[25]),  .B(n2977),  .C(n3088),  .D(b_reg[25]), .Y(n5535));
   NAND2X1 U6708 ( .A(digest[217]),  .B(n3045), .Y(n5534));
   OAI21X1 U6709 ( .A(n2126),  .B(n5536),  .C(n5537), .Y(puf_13_wire_3));
   AOI22X1 U6710 ( .A(a_reg[26]),  .B(n2977),  .C(digest[218]),  .D(n4718), .Y(n5537));
   NAND3X1 U6711 ( .A(n5538),  .B(n3090),  .C(n5539), .Y(n1335));
   AOI22X1 U6712 ( .A(a_reg[27]),  .B(n2979),  .C(n3088),  .D(b_reg[27]), .Y(n5539));
   NAND2X1 U6713 ( .A(digest[219]),  .B(n3045), .Y(n5538));
   NAND3X1 U6714 ( .A(n5540),  .B(n3091),  .C(n5541), .Y(n1334));
   AOI22X1 U6715 ( .A(a_reg[28]),  .B(n2977),  .C(b_reg[28]),  .D(n3088), .Y(n5541));
   NAND2X1 U6716 ( .A(digest[220]),  .B(n3045), .Y(n5540));
   NAND3X1 U6717 ( .A(n5542),  .B(n3090),  .C(n5543), .Y(n1333));
   AOI22X1 U6718 ( .A(a_reg[29]),  .B(n2978),  .C(n3089),  .D(b_reg[29]), .Y(n5543));
   NAND2X1 U6719 ( .A(digest[221]),  .B(n3045), .Y(n5542));
   OAI21X1 U6720 ( .A(n2126),  .B(n5544),  .C(n5545), .Y(n1332));
   AOI22X1 U6721 ( .A(a_reg[30]),  .B(n2977),  .C(digest[222]),  .D(n4718), .Y(n5545));
   NAND3X1 U6722 ( .A(n5546),  .B(n3090),  .C(n5547), .Y(n1331));
   AOI22X1 U6723 ( .A(a_reg[31]),  .B(n2977),  .C(b_reg[31]),  .D(n3088), .Y(n5547));
   NAND2X1 U6724 ( .A(digest[223]),  .B(n3045), .Y(n5546));
   OAI21X1 U6725 ( .A(n4713),  .B(n5548),  .C(n5549), .Y(n1330));
   AOI21X1 U6726 ( .A(N582),  .B(n3087),  .C(n4783), .Y(n5549));
   INVX1 U6727 ( .A(digest[192]), .Y(n5548));
   OAI21X1 U6728 ( .A(n3082),  .B(n5550),  .C(n2134), .Y(n1329));
   INVX1 U6729 ( .A(digest[193]), .Y(n5550));
   OAI21X1 U6730 ( .A(n3083),  .B(n5552),  .C(n2530), .Y(n1328));
   AOI21X1 U6731 ( .A(N584),  .B(n3087),  .C(n4783), .Y(n5553));
   INVX1 U6732 ( .A(digest[194]), .Y(n5552));
   OAI21X1 U6733 ( .A(n3082),  .B(n5554),  .C(n2144), .Y(n1327));
   INVX1 U6734 ( .A(digest[195]), .Y(n5554));
   OAI21X1 U6735 ( .A(n4713),  .B(n5556),  .C(n2157), .Y(n1326));
   INVX1 U6736 ( .A(digest[196]), .Y(n5556));
   OAI21X1 U6737 ( .A(n4713),  .B(n5558),  .C(n2269), .Y(n1325));
   INVX1 U6738 ( .A(digest[197]), .Y(n5558));
   OAI21X1 U6739 ( .A(n3083),  .B(n5560),  .C(n2319), .Y(n1324));
   INVX1 U6740 ( .A(digest[198]), .Y(n5560));
   OAI21X1 U6741 ( .A(n3083),  .B(n5562),  .C(n2191), .Y(n1323));
   AOI21X1 U6742 ( .A(N589),  .B(n3086),  .C(n4783), .Y(n5563));
   INVX1 U6743 ( .A(digest[199]), .Y(n5562));
   OAI21X1 U6744 ( .A(n3083),  .B(n5564),  .C(n2373), .Y(n1322));
   INVX1 U6745 ( .A(digest[200]), .Y(n5564));
   OAI21X1 U6746 ( .A(n3082),  .B(n5566),  .C(n2218), .Y(n1321));
   AOI21X1 U6747 ( .A(N591),  .B(n3085),  .C(n4783), .Y(n5567));
   INVX1 U6748 ( .A(digest[201]), .Y(n5566));
   OAI21X1 U6749 ( .A(n3083),  .B(n5568),  .C(n2261), .Y(n1320));
   AOI21X1 U6750 ( .A(N592),  .B(n3086),  .C(n4783), .Y(n5569));
   INVX1 U6751 ( .A(digest[202]), .Y(n5568));
   OAI21X1 U6752 ( .A(n4713),  .B(n5570),  .C(n2311), .Y(n1319));
   AOI21X1 U6753 ( .A(N593),  .B(n3085),  .C(n3093), .Y(n5571));
   INVX1 U6754 ( .A(digest[203]), .Y(n5570));
   OAI21X1 U6755 ( .A(n3083),  .B(n5572),  .C(n2176), .Y(n1318));
   INVX1 U6756 ( .A(digest[204]), .Y(n5572));
   OAI21X1 U6757 ( .A(n3083),  .B(n5574),  .C(n2365), .Y(n1317));
   AOI21X1 U6758 ( .A(N595),  .B(n3085),  .C(n4783), .Y(n5575));
   INVX1 U6759 ( .A(digest[205]), .Y(n5574));
   OAI21X1 U6760 ( .A(n3082),  .B(n5576),  .C(n2197), .Y(n1316));
   INVX1 U6761 ( .A(digest[206]), .Y(n5576));
   OAI21X1 U6762 ( .A(n4713),  .B(n5578),  .C(n2707), .Y(n1315));
   AOI21X1 U6763 ( .A(N597),  .B(n3085),  .C(n3093), .Y(n5579));
   INVX1 U6764 ( .A(digest[207]), .Y(n5578));
   OAI21X1 U6765 ( .A(n4713),  .B(n5580),  .C(n2421), .Y(n1314));
   AOI21X1 U6766 ( .A(N598),  .B(n3085),  .C(n4783), .Y(n5581));
   INVX1 U6767 ( .A(digest[208]), .Y(n5580));
   OAI21X1 U6768 ( .A(n4713),  .B(n5582),  .C(n2771), .Y(n1313));
   AOI21X1 U6769 ( .A(N599),  .B(n3085),  .C(n3093), .Y(n5583));
   INVX1 U6770 ( .A(digest[209]), .Y(n5582));
   OAI21X1 U6771 ( .A(n3082),  .B(n5584),  .C(n2834), .Y(n1312));
   AOI21X1 U6772 ( .A(N600),  .B(n3087),  .C(n4783), .Y(n5585));
   INVX1 U6773 ( .A(digest[210]), .Y(n5584));
   OAI21X1 U6774 ( .A(n3083),  .B(n5586),  .C(n2226), .Y(n1311));
   INVX1 U6775 ( .A(digest[211]), .Y(n5586));
   OAI21X1 U6776 ( .A(n4713),  .B(n5588),  .C(n2430), .Y(n1310));
   INVX1 U6777 ( .A(digest[212]), .Y(n5588));
   OAI21X1 U6778 ( .A(n4713),  .B(n5590),  .C(n2941), .Y(n1309));
   AOI21X1 U6779 ( .A(N603),  .B(n3085),  .C(n4783), .Y(n5591));
   INVX1 U6780 ( .A(digest[213]), .Y(n5590));
   OAI21X1 U6781 ( .A(n4713),  .B(n5592),  .C(n2170), .Y(n1308));
   AOI21X1 U6782 ( .A(N604),  .B(n3086),  .C(n3093), .Y(n5593));
   INVX1 U6783 ( .A(digest[214]), .Y(n5592));
   OAI21X1 U6784 ( .A(n3083),  .B(n5594),  .C(n2486), .Y(n1307));
   INVX1 U6785 ( .A(digest[215]), .Y(n5594));
   OAI21X1 U6786 ( .A(n3083),  .B(n5596),  .C(n2219), .Y(n1306));
   AOI21X1 U6787 ( .A(N606),  .B(n3087),  .C(n3093), .Y(n5597));
   INVX1 U6788 ( .A(digest[216]), .Y(n5596));
   OAI21X1 U6789 ( .A(n3082),  .B(n5598),  .C(n2312), .Y(n1305));
   AOI21X1 U6790 ( .A(N607),  .B(n3085),  .C(n4783), .Y(n5599));
   INVX1 U6791 ( .A(digest[217]), .Y(n5598));
   OAI21X1 U6792 ( .A(n3083),  .B(n5600),  .C(n2600), .Y(n1304));
   INVX1 U6793 ( .A(digest[218]), .Y(n5600));
   OAI21X1 U6794 ( .A(n3083),  .B(n5602),  .C(n2192), .Y(n1303));
   AOI21X1 U6795 ( .A(N609),  .B(n3086),  .C(n3093), .Y(n5603));
   INVX1 U6796 ( .A(digest[219]), .Y(n5602));
   OAI21X1 U6797 ( .A(n4713),  .B(n5604),  .C(n2366), .Y(n1302));
   AOI21X1 U6798 ( .A(N610),  .B(n3085),  .C(n3093), .Y(n5605));
   INVX1 U6799 ( .A(digest[220]), .Y(n5604));
   OAI21X1 U6800 ( .A(n3082),  .B(n5606),  .C(n2588), .Y(n1301));
   AOI21X1 U6801 ( .A(N611),  .B(n3086),  .C(n3093), .Y(n5607));
   INVX1 U6802 ( .A(digest[221]), .Y(n5606));
   OAI21X1 U6803 ( .A(n3083),  .B(n5608),  .C(n2662), .Y(n1300));
   INVX1 U6804 ( .A(digest[222]), .Y(n5608));
   OAI21X1 U6805 ( .A(n3083),  .B(n5610),  .C(n5611), .Y(n1299));
   AOI21X1 U6806 ( .A(N613),  .B(n3087),  .C(n3093), .Y(n5611));
   INVX1 U6807 ( .A(digest[223]), .Y(n5610));
   OAI21X1 U6808 ( .A(n2126),  .B(n5612),  .C(n5613), .Y(n1298));
   AOI22X1 U6809 ( .A(b_reg[0]),  .B(n2979),  .C(digest[160]),  .D(n4718), .Y(n5613));
   INVX1 U6810 ( .A(c_reg[0]), .Y(n5612));
   NAND3X1 U6811 ( .A(n5614),  .B(n3090),  .C(n5615), .Y(n1297));
   AOI22X1 U6812 ( .A(b_reg[1]),  .B(n2978),  .C(c_reg[1]),  .D(n3089), .Y(n5615));
   NAND2X1 U6813 ( .A(digest[161]),  .B(n3045), .Y(n5614));
   OAI21X1 U6814 ( .A(n5616),  .B(n2126),  .C(n5617), .Y(n1296));
   AOI22X1 U6815 ( .A(b_reg[2]),  .B(n2977),  .C(digest[162]),  .D(n4718), .Y(n5617));
   INVX1 U6816 ( .A(c_reg[2]), .Y(n5616));
   OAI21X1 U6817 ( .A(n2126),  .B(n5618),  .C(n5619), .Y(n1295));
   AOI22X1 U6818 ( .A(b_reg[3]),  .B(n2979),  .C(digest[163]),  .D(n4718), .Y(n5619));
   INVX1 U6819 ( .A(c_reg[3]), .Y(n5618));
   NAND3X1 U6820 ( .A(n5620),  .B(n3090),  .C(n5621), .Y(n1294));
   AOI22X1 U6821 ( .A(b_reg[4]),  .B(n2977),  .C(c_reg[4]),  .D(n3088), .Y(n5621));
   NAND2X1 U6822 ( .A(digest[164]),  .B(n3045), .Y(puf_14_wire_3));
   NAND3X1 U6823 ( .A(n5622),  .B(n3090),  .C(n5623), .Y(n1293));
   AOI22X1 U6824 ( .A(b_reg[5]),  .B(n2977),  .C(c_reg[5]),  .D(n3089), .Y(n5623));
   NAND2X1 U6825 ( .A(digest[165]),  .B(n3045), .Y(n5622));
   NAND3X1 U6826 ( .A(n5624),  .B(n3091),  .C(n5625), .Y(n1292));
   AOI22X1 U6827 ( .A(b_reg[6]),  .B(n2979),  .C(c_reg[6]),  .D(n3089), .Y(n5625));
   NAND2X1 U6828 ( .A(digest[166]),  .B(n3045), .Y(n5624));
   OAI21X1 U6829 ( .A(n2126),  .B(n5626),  .C(n5627), .Y(n1291));
   AOI22X1 U6830 ( .A(b_reg[7]),  .B(n2980),  .C(digest[167]),  .D(n4718), .Y(n5627));
   INVX1 U6831 ( .A(c_reg[7]), .Y(n5626));
   NAND3X1 U6832 ( .A(n5628),  .B(n3090),  .C(n5629), .Y(n1290));
   AOI22X1 U6833 ( .A(b_reg[8]),  .B(n2977),  .C(c_reg[8]),  .D(n3089), .Y(n5629));
   NAND2X1 U6834 ( .A(digest[168]),  .B(n3045), .Y(n5628));
   NAND3X1 U6835 ( .A(n5630),  .B(n3090),  .C(n5631), .Y(n1289));
   AOI22X1 U6836 ( .A(b_reg[9]),  .B(n2980),  .C(n3089),  .D(c_reg[9]), .Y(n5631));
   NAND2X1 U6837 ( .A(digest[169]),  .B(n3045), .Y(n5630));
   OAI21X1 U6838 ( .A(n5632),  .B(n2126),  .C(n5633), .Y(n1288));
   AOI22X1 U6839 ( .A(b_reg[10]),  .B(n2977),  .C(digest[170]),  .D(n4718), .Y(n5633));
   INVX1 U6840 ( .A(c_reg[10]), .Y(n5632));
   OAI21X1 U6841 ( .A(n2126),  .B(n5634),  .C(n5635), .Y(n1287));
   AOI22X1 U6842 ( .A(b_reg[11]),  .B(n2979),  .C(digest[171]),  .D(n4718), .Y(n5635));
   INVX1 U6843 ( .A(c_reg[11]), .Y(n5634));
   NAND3X1 U6844 ( .A(n5636),  .B(n3091),  .C(n5637), .Y(n1286));
   AOI22X1 U6845 ( .A(b_reg[12]),  .B(n2979),  .C(c_reg[12]),  .D(n3089), .Y(n5637));
   NAND2X1 U6846 ( .A(digest[172]),  .B(n3045), .Y(n5636));
   NAND3X1 U6847 ( .A(n5638),  .B(n3091),  .C(n5639), .Y(n1285));
   AOI22X1 U6848 ( .A(b_reg[13]),  .B(n2978),  .C(c_reg[13]),  .D(n3089), .Y(n5639));
   NAND2X1 U6849 ( .A(digest[173]),  .B(n3045), .Y(n5638));
   NAND3X1 U6850 ( .A(n5640),  .B(n3091),  .C(n5641), .Y(n1284));
   AOI22X1 U6851 ( .A(b_reg[14]),  .B(n2977),  .C(c_reg[14]),  .D(n3089), .Y(n5641));
   NAND2X1 U6852 ( .A(digest[174]),  .B(n3045), .Y(n5640));
   NAND3X1 U6853 ( .A(n5642),  .B(n3090),  .C(n1909), .Y(n1283));
   AOI22X1 U6854 ( .A(b_reg[15]),  .B(n2978),  .C(c_reg[15]),  .D(n3089), .Y(n5643));
   NAND2X1 U6855 ( .A(digest[175]),  .B(n3045), .Y(n5642));
   OAI21X1 U6856 ( .A(n2126),  .B(n5644),  .C(n5645), .Y(n1282));
   AOI22X1 U6857 ( .A(b_reg[16]),  .B(n2979),  .C(digest[176]),  .D(n4718), .Y(n5645));
   INVX1 U6858 ( .A(c_reg[16]), .Y(n5644));
   NAND3X1 U6859 ( .A(n5646),  .B(n3090),  .C(n1910), .Y(n1281));
   AOI22X1 U6860 ( .A(b_reg[17]),  .B(n2980),  .C(c_reg[17]),  .D(n3089), .Y(n5647));
   NAND2X1 U6861 ( .A(digest[177]),  .B(n3045), .Y(n5646));
   NAND3X1 U6862 ( .A(n5648),  .B(n3091),  .C(n1911), .Y(n1280));
   AOI22X1 U6863 ( .A(b_reg[18]),  .B(n2978),  .C(c_reg[18]),  .D(n3089), .Y(n5649));
   NAND2X1 U6864 ( .A(digest[178]),  .B(n3045), .Y(n5648));
   NAND3X1 U6865 ( .A(n5650),  .B(n3091),  .C(n1912), .Y(n1279));
   AOI22X1 U6866 ( .A(b_reg[19]),  .B(n2980),  .C(c_reg[19]),  .D(n3089), .Y(n5651));
   NAND2X1 U6867 ( .A(digest[179]),  .B(n3046), .Y(n5650));
   OAI21X1 U6868 ( .A(n2126),  .B(n5652),  .C(n5653), .Y(n1278));
   AOI22X1 U6869 ( .A(b_reg[20]),  .B(n2978),  .C(digest[180]),  .D(n4718), .Y(n5653));
   INVX1 U6870 ( .A(c_reg[20]), .Y(n5652));
   NAND3X1 U6871 ( .A(n5654),  .B(n3090),  .C(n1913), .Y(n1277));
   AOI22X1 U6872 ( .A(b_reg[21]),  .B(n2980),  .C(c_reg[21]),  .D(n3089), .Y(n5655));
   NAND2X1 U6873 ( .A(digest[181]),  .B(n3046), .Y(n5654));
   NAND3X1 U6874 ( .A(n5656),  .B(n3091),  .C(n1914), .Y(n1276));
   AOI22X1 U6875 ( .A(b_reg[22]),  .B(n2977),  .C(c_reg[22]),  .D(n3089), .Y(n5657));
   NAND2X1 U6876 ( .A(digest[182]),  .B(n3046), .Y(n5656));
   OAI21X1 U6877 ( .A(n2126),  .B(n5658),  .C(n5659), .Y(n1275));
   AOI22X1 U6878 ( .A(b_reg[23]),  .B(n2979),  .C(digest[183]),  .D(n4718), .Y(n5659));
   INVX1 U6879 ( .A(c_reg[23]), .Y(n5658));
   OAI21X1 U6880 ( .A(n2126),  .B(n5660),  .C(n5661), .Y(n1274));
   AOI22X1 U6881 ( .A(b_reg[24]),  .B(n2978),  .C(digest[184]),  .D(n4718), .Y(n5661));
   INVX1 U6882 ( .A(c_reg[24]), .Y(n5660));
   OAI21X1 U6883 ( .A(n5662),  .B(n2126),  .C(n5663), .Y(n1273));
   AOI22X1 U6884 ( .A(b_reg[25]),  .B(n2977),  .C(digest[185]),  .D(n4718), .Y(n5663));
   INVX1 U6885 ( .A(c_reg[25]), .Y(n5662));
   NAND3X1 U6886 ( .A(n5664),  .B(n3091),  .C(n1915), .Y(n1272));
   AOI22X1 U6887 ( .A(b_reg[26]),  .B(n2979),  .C(c_reg[26]),  .D(n3089), .Y(n5665));
   NAND2X1 U6888 ( .A(digest[186]),  .B(n3046), .Y(n5664));
   NAND3X1 U6889 ( .A(n5666),  .B(n3091),  .C(n1916), .Y(n1271));
   AOI22X1 U6890 ( .A(b_reg[27]),  .B(n2978),  .C(n3089),  .D(c_reg[27]), .Y(n5667));
   NAND2X1 U6891 ( .A(digest[187]),  .B(n3046), .Y(n5666));
   NAND3X1 U6892 ( .A(n5668),  .B(n3091),  .C(n1917), .Y(n1270));
   AOI22X1 U6893 ( .A(b_reg[28]),  .B(n2980),  .C(c_reg[28]),  .D(n3088), .Y(n5669));
   NAND2X1 U6894 ( .A(digest[188]),  .B(n3046), .Y(n5668));
   NAND3X1 U6895 ( .A(n5670),  .B(n3090),  .C(n1918), .Y(n1269));
   AOI22X1 U6896 ( .A(b_reg[29]),  .B(n2979),  .C(n3089),  .D(c_reg[29]), .Y(n5671));
   NAND2X1 U6897 ( .A(digest[189]),  .B(n3046), .Y(n5670));
   OAI21X1 U6898 ( .A(n2126),  .B(n5672),  .C(n5673), .Y(n1268));
   AOI22X1 U6899 ( .A(b_reg[30]),  .B(n2979),  .C(digest[190]),  .D(n4718), .Y(n5673));
   INVX1 U6900 ( .A(c_reg[30]), .Y(n5672));
   OAI21X1 U6901 ( .A(n2126),  .B(n5674),  .C(n5675), .Y(n1267));
   AOI22X1 U6902 ( .A(b_reg[31]),  .B(n2977),  .C(digest[191]),  .D(n4718), .Y(n5675));
   NAND3X1 U6903 ( .A(n3100),  .B(n4692),  .C(sha256_ctrl_reg[0]), .Y(n4699));
   INVX1 U6904 ( .A(c_reg[31]), .Y(n5674));
   OAI21X1 U6905 ( .A(next),  .B(init),  .C(ready), .Y(n3116));
   AND2X1 U6906 ( .A(n4695),  .B(n4692), .Y(ready));
   INVX1 U6907 ( .A(sha256_ctrl_reg[1]), .Y(n4692));
   OAI21X1 U6908 ( .A(n4713),  .B(n5677),  .C(n2725), .Y(n1266));
   INVX1 U6909 ( .A(digest[160]), .Y(n5677));
   OAI21X1 U6910 ( .A(n3082),  .B(n5679),  .C(n2476), .Y(n1265));
   AOI21X1 U6911 ( .A(N615),  .B(n3087),  .C(n3093), .Y(n5680));
   INVX1 U6912 ( .A(digest[161]), .Y(n5679));
   OAI21X1 U6913 ( .A(n4713),  .B(n5681),  .C(n2788), .Y(n1264));
   INVX1 U6914 ( .A(digest[162]), .Y(n5681));
   OAI21X1 U6915 ( .A(n3083),  .B(n5683),  .C(n2544), .Y(n1263));
   INVX1 U6916 ( .A(digest[163]), .Y(n5683));
   OAI21X1 U6917 ( .A(n3083),  .B(n5685),  .C(n2645), .Y(n1262));
   AOI21X1 U6918 ( .A(N618),  .B(n3086),  .C(n4783), .Y(n5686));
   INVX1 U6919 ( .A(digest[164]), .Y(n5685));
   OAI21X1 U6920 ( .A(n3082),  .B(n5687),  .C(n2708), .Y(n1261));
   AOI21X1 U6921 ( .A(N619),  .B(n3087),  .C(n3093), .Y(n5688));
   INVX1 U6922 ( .A(digest[165]), .Y(n5687));
   OAI21X1 U6923 ( .A(n3082),  .B(n5689),  .C(n2835), .Y(n1260));
   AOI21X1 U6924 ( .A(N620),  .B(n3085),  .C(n4783), .Y(n5690));
   INVX1 U6925 ( .A(digest[166]), .Y(n5689));
   OAI21X1 U6926 ( .A(n3083),  .B(n5691),  .C(n2320), .Y(n1259));
   INVX1 U6927 ( .A(digest[167]), .Y(n5691));
   OAI21X1 U6928 ( .A(n3083),  .B(n5693),  .C(n2772), .Y(n1258));
   AOI21X1 U6929 ( .A(N622),  .B(n3086),  .C(n4783), .Y(n5694));
   INVX1 U6930 ( .A(digest[168]), .Y(n5693));
   OAI21X1 U6931 ( .A(n3082),  .B(n5695),  .C(n2942), .Y(n1257));
   AOI21X1 U6932 ( .A(N623),  .B(n3086),  .C(n4783), .Y(n5696));
   INVX1 U6933 ( .A(digest[169]), .Y(n5695));
   OAI21X1 U6934 ( .A(n3082),  .B(n5697),  .C(n2374), .Y(n1256));
   INVX1 U6935 ( .A(digest[170]), .Y(n5697));
   OAI21X1 U6936 ( .A(n3082),  .B(n5699),  .C(n2487), .Y(n1255));
   INVX1 U6937 ( .A(digest[171]), .Y(n5699));
   OAI21X1 U6938 ( .A(n4713),  .B(n5701),  .C(n2262), .Y(n1254));
   AOI21X1 U6939 ( .A(N626),  .B(n3087),  .C(n4783), .Y(n5702));
   INVX1 U6940 ( .A(digest[172]), .Y(n5701));
   OAI21X1 U6941 ( .A(n3082),  .B(n5703),  .C(n2220), .Y(n1253));
   AOI21X1 U6942 ( .A(N627),  .B(n3086),  .C(n4783), .Y(n5704));
   INVX1 U6943 ( .A(digest[173]), .Y(n5703));
   OAI21X1 U6944 ( .A(n3082),  .B(n5705),  .C(n2313), .Y(n1252));
   AOI21X1 U6945 ( .A(N628),  .B(n3086),  .C(n4783), .Y(n5706));
   INVX1 U6946 ( .A(digest[174]), .Y(n5705));
   OAI21X1 U6947 ( .A(n3082),  .B(n5707),  .C(n2367), .Y(n1251));
   AOI21X1 U6948 ( .A(N629),  .B(n3086),  .C(n4783), .Y(n5708));
   INVX1 U6949 ( .A(digest[175]), .Y(n5707));
   OAI21X1 U6950 ( .A(n3082),  .B(n5709),  .C(n2227), .Y(n1250));
   INVX1 U6951 ( .A(digest[176]), .Y(n5709));
   OAI21X1 U6952 ( .A(n3083),  .B(n5711),  .C(n2422), .Y(n1249));
   AOI21X1 U6953 ( .A(N631),  .B(n3085),  .C(n4783), .Y(n5712));
   INVX1 U6954 ( .A(digest[177]), .Y(n5711));
   OAI21X1 U6955 ( .A(n3083),  .B(n5713),  .C(n2531), .Y(n1248));
   AOI21X1 U6956 ( .A(N632),  .B(n3087),  .C(n4783), .Y(n5714));
   INVX1 U6957 ( .A(digest[178]), .Y(n5713));
   OAI21X1 U6958 ( .A(n3082),  .B(n5715),  .C(n2646), .Y(n1247));
   AOI21X1 U6959 ( .A(N633),  .B(n3086),  .C(n4783), .Y(n5716));
   INVX1 U6960 ( .A(digest[179]), .Y(n5715));
   OAI21X1 U6961 ( .A(n3083),  .B(n5717),  .C(n2270), .Y(n1246));
   INVX1 U6962 ( .A(digest[180]), .Y(n5717));
   OAI21X1 U6963 ( .A(n4713),  .B(n5719),  .C(n2773), .Y(n1245));
   AOI21X1 U6964 ( .A(N635),  .B(n3087),  .C(n4783), .Y(n5720));
   INVX1 U6965 ( .A(digest[181]), .Y(n5719));
   OAI21X1 U6966 ( .A(n4713),  .B(n5721),  .C(n2709), .Y(n1244));
   AOI21X1 U6967 ( .A(N636),  .B(n3086),  .C(n3093), .Y(n5722));
   INVX1 U6968 ( .A(digest[182]), .Y(n5721));
   OAI21X1 U6969 ( .A(n3083),  .B(n5723),  .C(n2431), .Y(n1243));
   INVX1 U6970 ( .A(digest[183]), .Y(n5723));
   OAI21X1 U6971 ( .A(n3082),  .B(n5725),  .C(n2545), .Y(n1242));
   INVX1 U6972 ( .A(digest[184]), .Y(n5725));
   OAI21X1 U6973 ( .A(n4713),  .B(n5727),  .C(n2898), .Y(n1241));
   INVX1 U6974 ( .A(digest[185]), .Y(n5727));
   OAI21X1 U6975 ( .A(n3082),  .B(n5729),  .C(n2836), .Y(n1240));
   AOI21X1 U6976 ( .A(N640),  .B(n3087),  .C(n4783), .Y(n5730));
   INVX1 U6977 ( .A(digest[186]), .Y(n5729));
   OAI21X1 U6978 ( .A(n3083),  .B(n5731),  .C(n2477), .Y(n1239));
   AOI21X1 U6979 ( .A(N641),  .B(n3087),  .C(n3093), .Y(n5732));
   INVX1 U6980 ( .A(digest[187]), .Y(n5731));
   OAI21X1 U6981 ( .A(n3083),  .B(n5733),  .C(n2589), .Y(n1238));
   AOI21X1 U6982 ( .A(N642),  .B(n3086),  .C(n3093), .Y(n5734));
   INVX1 U6983 ( .A(digest[188]), .Y(n5733));
   OAI21X1 U6984 ( .A(n3082),  .B(n5735),  .C(n2943), .Y(n1237));
   AOI21X1 U6985 ( .A(N643),  .B(n3086),  .C(n3093), .Y(n5736));
   INVX1 U6986 ( .A(digest[189]), .Y(n5735));
   OAI21X1 U6987 ( .A(n3083),  .B(n5738),  .C(n2789), .Y(n1236));
   INVX1 U6988 ( .A(digest[190]), .Y(n5738));
   OAI21X1 U6989 ( .A(n3083),  .B(n5740),  .C(n2949), .Y(n1235));
   NAND3X1 U6990 ( .A(n3100),  .B(n4695),  .C(sha256_ctrl_reg[1]), .Y(n4696));
   INVX1 U6991 ( .A(rst), .Y(n3100));
   INVX1 U6992 ( .A(digest[191]), .Y(n5740));
   OAI21X1 U6993 ( .A(sha256_ctrl_reg[0]),  .B(n5676),  .C(n2951), .Y(n4713));
   AOI21X1 U6994 ( .A(n4695),  .B(sha256_ctrl_reg[1]),  .C(rst), .Y(n5737));
   INVX1 U6995 ( .A(sha256_ctrl_reg[0]), .Y(n4695));
   INVX1 U6996 ( .A(init), .Y(n5676));
   INVX1 U6997 ( .A(n5745), .Y(n5744));
   NAND3X1 U6998 ( .A(n5746),  .B(n5747),  .C(n5748), .Y(n5745));
   OAI21X1 U6999 ( .A(n2846),  .B(n1978),  .C(n5917), .Y(n5748));
   NAND3X1 U7000 ( .A(n6000),  .B(n4705),  .C(n2893), .Y(n5747));
   NOR3X1 U7001 ( .A(n6050),  .B(n5752),  .C(n6069), .Y(n5746));
   AOI22X1 U7002 ( .A(n5789),  .B(n5753),  .C(n6061),  .D(n2656), .Y(n5743));
   OR2X1 U7003 ( .A(n2110),  .B(n1973), .Y(n5753));
   AOI22X1 U7004 ( .A(n5860),  .B(n6001),  .C(n5763),  .D(n2717), .Y(n5742));
   AOI21X1 U7005 ( .A(n5917),  .B(n5760),  .C(n5761), .Y(n5759));
   OAI21X1 U7006 ( .A(n5762),  .B(n2720),  .C(n5764), .Y(n5761));
   OAI21X1 U7007 ( .A(n5972),  .B(n2846),  .C(n5789), .Y(n5764));
   AND2X1 U7008 ( .A(n5765),  .B(n5766), .Y(n5762));
   AOI22X1 U7009 ( .A(n5859),  .B(n6021),  .C(n5846),  .D(n4707), .Y(n5766));
   AOI21X1 U7010 ( .A(n5934),  .B(t_ctr_reg[5]),  .C(n5767), .Y(n5765));
   NAND3X1 U7011 ( .A(n5768),  .B(n2114),  .C(n5770), .Y(n5760));
   INVX1 U7012 ( .A(n1965), .Y(n5768));
   AOI21X1 U7013 ( .A(n5934),  .B(n6001),  .C(n5774), .Y(n5758));
   INVX1 U7014 ( .A(n5775), .Y(k_data[7]));
   NOR3X1 U7015 ( .A(n1775),  .B(n1945),  .C(n1948), .Y(n5775));
   NAND3X1 U7016 ( .A(n2112),  .B(n2109),  .C(n1930), .Y(n5777));
   NAND3X1 U7017 ( .A(n2101),  .B(n2892),  .C(n1966), .Y(n5776));
   AOI21X1 U7018 ( .A(n5904),  .B(n2956),  .C(n5787), .Y(n5785));
   OAI21X1 U7019 ( .A(n1957),  .B(n2849),  .C(n5790), .Y(n5787));
   OAI21X1 U7020 ( .A(n5821),  .B(n1977),  .C(n6001), .Y(n5790));
   AOI22X1 U7021 ( .A(n5917),  .B(n2652),  .C(n5846),  .D(n2848), .Y(n5784));
   OR2X1 U7022 ( .A(n5794),  .B(n5795), .Y(k_data[6]));
   NAND3X1 U7023 ( .A(n5796),  .B(n5797),  .C(n1919), .Y(n5795));
   AOI22X1 U7024 ( .A(n6001),  .B(n1972),  .C(n5885),  .D(n5763), .Y(n5798));
   INVX1 U7025 ( .A(n5800), .Y(n5797));
   INVX1 U7026 ( .A(n1954), .Y(n5796));
   NAND3X1 U7027 ( .A(n5802),  .B(n1962),  .C(n1920), .Y(n5794));
   AOI22X1 U7028 ( .A(n5789),  .B(n5805),  .C(n5981),  .D(t_ctr_reg[2]), .Y(n5804));
   NAND2X1 U7029 ( .A(n5917),  .B(n5806), .Y(n5802));
   OAI21X1 U7030 ( .A(t_ctr_reg[4]),  .B(n2593),  .C(n2892), .Y(n5806));
   NOR3X1 U7031 ( .A(n5811),  .B(n1976),  .C(n5813), .Y(n5810));
   OAI21X1 U7032 ( .A(n5848),  .B(n2953),  .C(n5815), .Y(n5811));
   AOI22X1 U7033 ( .A(n5874),  .B(n2785),  .C(n5845),  .D(n2893), .Y(n5815));
   AOI21X1 U7034 ( .A(n5789),  .B(n5998),  .C(n5817), .Y(n5809));
   NAND2X1 U7035 ( .A(n5818),  .B(n2653), .Y(n5817));
   OAI21X1 U7036 ( .A(n5831),  .B(n1963),  .C(n5763), .Y(n5818));
   AOI22X1 U7037 ( .A(n6001),  .B(n1978),  .C(n5772),  .D(n5917), .Y(n5808));
   NOR3X1 U7038 ( .A(n5826),  .B(n5752),  .C(n5783), .Y(n5825));
   OAI21X1 U7039 ( .A(n2424),  .B(n2849),  .C(n5828), .Y(n5826));
   OAI21X1 U7040 ( .A(n5821),  .B(n5845),  .C(n2785), .Y(n5828));
   AOI21X1 U7041 ( .A(t_ctr_reg[3]),  .B(n4711),  .C(n5859), .Y(n5827));
   AOI22X1 U7042 ( .A(n5917),  .B(n5829),  .C(n6001),  .D(n1980), .Y(n5824));
   NAND3X1 U7043 ( .A(n2783),  .B(n2889),  .C(n5832), .Y(n5829));
   AOI22X1 U7044 ( .A(n5814),  .B(n2893),  .C(n5934),  .D(n5763), .Y(n5823));
   INVX1 U7045 ( .A(n5836), .Y(n5835));
   NAND3X1 U7046 ( .A(n5837),  .B(n2653),  .C(n2111), .Y(n5836));
   OAI21X1 U7047 ( .A(n5904),  .B(n5934),  .C(n5917), .Y(n5839));
   AOI22X1 U7048 ( .A(n5789),  .B(n5841),  .C(n6001),  .D(n5842), .Y(n5834));
   NAND3X1 U7049 ( .A(n2842),  .B(n2892),  .C(n1931), .Y(n5842));
   OR2X1 U7050 ( .A(n1972),  .B(n2110), .Y(n5841));
   AOI22X1 U7051 ( .A(n1981),  .B(n2784),  .C(n5763),  .D(n2716), .Y(n5833));
   NOR3X1 U7052 ( .A(n2535),  .B(n5853),  .C(n5854), .Y(n5851));
   OAI21X1 U7053 ( .A(n5822),  .B(n2846),  .C(n5763), .Y(n5856));
   OAI21X1 U7054 ( .A(n5857),  .B(n5858),  .C(n2956), .Y(n5855));
   OAI21X1 U7055 ( .A(n6021),  .B(n2594),  .C(n2654), .Y(n5858));
   NAND3X1 U7056 ( .A(n2889),  .B(n2847),  .C(n2593), .Y(n5857));
   AOI22X1 U7057 ( .A(n5772),  .B(n5789),  .C(n5936),  .D(n2955), .Y(n5850));
   OR2X1 U7058 ( .A(n5862),  .B(n5863), .Y(k_data[30]));
   NAND3X1 U7059 ( .A(n5864),  .B(n1961),  .C(n1921), .Y(n5863));
   AOI22X1 U7060 ( .A(n5867),  .B(n2955),  .C(n5925),  .D(n2848), .Y(n5866));
   INVX1 U7061 ( .A(n5868), .Y(n5864));
   NAND3X1 U7062 ( .A(n5869),  .B(n5870),  .C(n1922), .Y(n5862));
   AOI22X1 U7063 ( .A(n5789),  .B(n5872),  .C(n5873),  .D(n4703), .Y(n5871));
   NAND2X1 U7064 ( .A(n2890),  .B(n2655), .Y(n5872));
   NAND3X1 U7065 ( .A(t_ctr_reg[3]),  .B(n4707),  .C(n5886), .Y(n5870));
   NOR2X1 U7066 ( .A(n5752),  .B(n5981), .Y(n5869));
   NOR3X1 U7067 ( .A(n1937),  .B(n5880),  .C(n5881), .Y(n5878));
   INVX1 U7068 ( .A(n5882), .Y(n5881));
   OAI21X1 U7069 ( .A(n5771),  .B(n5821),  .C(n2656), .Y(n5882));
   NAND3X1 U7070 ( .A(n2101),  .B(n2104),  .C(n2111), .Y(n5879));
   AOI21X1 U7071 ( .A(n5782),  .B(n2848),  .C(n5884), .Y(n5877));
   OAI21X1 U7072 ( .A(n2844),  .B(n2103),  .C(n5887), .Y(n5884));
   NAND2X1 U7073 ( .A(n5789),  .B(n5888), .Y(n5887));
   NAND3X1 U7074 ( .A(n2114),  .B(n2115),  .C(n1932), .Y(n5888));
   AOI21X1 U7075 ( .A(n5874),  .B(n2893),  .C(n5891), .Y(n5876));
   OR2X1 U7076 ( .A(n5892),  .B(n5893), .Y(k_data[29]));
   NAND3X1 U7077 ( .A(n5894),  .B(n5895),  .C(n5896), .Y(n5893));
   AND2X1 U7078 ( .A(n5897),  .B(n5898), .Y(n5896));
   AOI22X1 U7079 ( .A(n5789),  .B(n6109),  .C(n5821),  .D(n2956), .Y(n5897));
   NAND2X1 U7080 ( .A(n5925),  .B(n2785), .Y(n5895));
   AOI22X1 U7081 ( .A(n5782),  .B(n2592),  .C(n5918),  .D(n6001), .Y(n5894));
   NAND3X1 U7082 ( .A(n5900),  .B(n5901),  .C(n5902), .Y(n5892));
   NOR3X1 U7083 ( .A(n6067),  .B(n5752),  .C(n5883), .Y(n5902));
   NAND2X1 U7084 ( .A(n5807),  .B(n2955), .Y(n5901));
   AOI22X1 U7085 ( .A(n5763),  .B(n2713),  .C(n5917),  .D(n1965), .Y(n5900));
   NAND3X1 U7086 ( .A(n2655),  .B(n2954),  .C(n2106), .Y(n5773));
   INVX1 U7087 ( .A(n5910), .Y(n5909));
   NAND3X1 U7088 ( .A(n5911),  .B(n2954),  .C(n2780), .Y(n5910));
   OAI21X1 U7089 ( .A(n5767),  .B(n5875),  .C(n5763), .Y(n5911));
   AOI22X1 U7090 ( .A(n6001),  .B(n5913),  .C(n5904),  .D(n2785), .Y(n5908));
   NAND2X1 U7091 ( .A(n2113),  .B(n2115), .Y(n5913));
   AOI22X1 U7092 ( .A(n1960),  .B(n2719),  .C(n5821),  .D(n2592), .Y(n5906));
   AOI21X1 U7093 ( .A(n6061),  .B(n2784),  .C(n5800), .Y(n5905));
   OAI21X1 U7094 ( .A(n2891),  .B(n2843),  .C(n5919), .Y(n5800));
   AOI21X1 U7095 ( .A(n5860),  .B(n5789),  .C(n5880), .Y(n5919));
   NOR3X1 U7096 ( .A(n5923),  .B(n5883),  .C(n5854), .Y(n5922));
   AND2X1 U7097 ( .A(n5904),  .B(n5789), .Y(n5854));
   OAI21X1 U7098 ( .A(n5926),  .B(n2891),  .C(n5924), .Y(n5923));
   OAI21X1 U7099 ( .A(n5846),  .B(n1981),  .C(n2955), .Y(n5924));
   AOI22X1 U7100 ( .A(n5860),  .B(n2893),  .C(n5813),  .D(n4705), .Y(n5921));
   AOI21X1 U7101 ( .A(n6109),  .B(n5763),  .C(n5927), .Y(n5920));
   NAND3X1 U7102 ( .A(n2481),  .B(n5929),  .C(n5930), .Y(k_data[26]));
   AOI21X1 U7103 ( .A(n5917),  .B(n5875),  .C(n5891), .Y(n5932));
   OAI21X1 U7104 ( .A(n5848),  .B(n2954),  .C(n5933), .Y(n5891));
   AOI22X1 U7105 ( .A(n5917),  .B(n2713),  .C(n5843),  .D(n5789), .Y(n5933));
   INVX1 U7106 ( .A(n5935), .Y(n5931));
   OAI21X1 U7107 ( .A(n2720),  .B(n2595),  .C(n5937), .Y(n5935));
   AOI22X1 U7108 ( .A(n5914),  .B(n2656),  .C(n5821),  .D(n2848), .Y(n5937));
   NOR3X1 U7109 ( .A(n5803),  .B(n5782),  .C(n5752), .Y(n5929));
   AOI21X1 U7110 ( .A(n6001),  .B(n1979),  .C(n5939), .Y(n5928));
   NOR3X1 U7111 ( .A(n2781),  .B(n5861),  .C(n4711), .Y(n5939));
   NAND3X1 U7112 ( .A(n2538),  .B(n5941),  .C(n5942), .Y(k_data[25]));
   AOI22X1 U7113 ( .A(n5918),  .B(n6001),  .C(n6109),  .D(n2785), .Y(n5944));
   AOI21X1 U7114 ( .A(n5934),  .B(n5789),  .C(n5945), .Y(n5943));
   NOR3X1 U7115 ( .A(n1938),  .B(n5912),  .C(n5947), .Y(n5941));
   INVX1 U7116 ( .A(n5948), .Y(n5947));
   OAI21X1 U7117 ( .A(n1980),  .B(n5845),  .C(n5763), .Y(n5948));
   AOI21X1 U7118 ( .A(n5915),  .B(n2595),  .C(n2891), .Y(n5946));
   AOI22X1 U7119 ( .A(n1959),  .B(n2784),  .C(t_ctr_reg[3]),  .D(n5813), .Y(n5940));
   NOR3X1 U7120 ( .A(n1851),  .B(n5927),  .C(n5953), .Y(n5952));
   OAI21X1 U7121 ( .A(n5848),  .B(n2892),  .C(n5954), .Y(n5927));
   NAND3X1 U7122 ( .A(n5917),  .B(n4707),  .C(n5874), .Y(n5954));
   AOI21X1 U7123 ( .A(n6002),  .B(t_ctr_reg[4]),  .C(n5981), .Y(n5951));
   AOI22X1 U7124 ( .A(n5889),  .B(n5789),  .C(n5821),  .D(n2719), .Y(n5950));
   NAND3X1 U7125 ( .A(n5955),  .B(n5956),  .C(n5957), .Y(k_data[23]));
   NOR3X1 U7126 ( .A(n5958),  .B(n5959),  .C(n1969), .Y(n5957));
   OAI21X1 U7127 ( .A(n5861),  .B(n2890),  .C(n5961), .Y(n5958));
   AOI22X1 U7128 ( .A(n5972),  .B(n2956),  .C(n5789),  .D(n1973), .Y(n5961));
   NOR3X1 U7129 ( .A(n5962),  .B(n5843),  .C(n5853), .Y(n5956));
   INVX1 U7130 ( .A(n2479), .Y(n5962));
   AOI21X1 U7131 ( .A(n5917),  .B(n5998),  .C(n5964), .Y(n5955));
   NAND2X1 U7132 ( .A(n5965),  .B(n2109), .Y(n5964));
   NAND3X1 U7133 ( .A(n5763),  .B(t_ctr_reg[5]),  .C(n5925), .Y(n5965));
   AOI21X1 U7134 ( .A(n5917),  .B(n5970),  .C(n6003), .Y(n5969));
   NAND2X1 U7135 ( .A(n5971),  .B(n2714), .Y(n5970));
   AOI22X1 U7136 ( .A(n6001),  .B(n5973),  .C(n5763),  .D(n2108), .Y(n5968));
   NAND3X1 U7137 ( .A(n2889),  .B(n2954),  .C(n2654), .Y(n5973));
   NAND3X1 U7138 ( .A(n5974),  .B(n2112),  .C(n1923), .Y(n5960));
   AOI22X1 U7139 ( .A(n5925),  .B(n5886),  .C(n5914),  .D(n5789), .Y(n5975));
   OAI21X1 U7140 ( .A(n5874),  .B(n5782),  .C(n5917), .Y(n5974));
   AOI22X1 U7141 ( .A(n5807),  .B(n2956),  .C(n5771),  .D(n2848), .Y(n5966));
   NOR3X1 U7142 ( .A(n5979),  .B(n1756),  .C(n5980), .Y(n5978));
   OAI21X1 U7143 ( .A(n2720),  .B(n2892),  .C(n5982), .Y(n5979));
   AOI22X1 U7144 ( .A(n5914),  .B(n2955),  .C(n6109),  .D(n2785), .Y(n5982));
   AOI21X1 U7145 ( .A(n5781),  .B(n6021),  .C(n5983), .Y(n5977));
   OAI21X1 U7146 ( .A(n5820),  .B(n2891),  .C(n5984), .Y(n5983));
   OAI21X1 U7147 ( .A(n5998),  .B(n2652),  .C(n6001), .Y(n5984));
   AOI22X1 U7148 ( .A(n5821),  .B(n2592),  .C(n5789),  .D(n2846), .Y(n5976));
   NAND3X1 U7149 ( .A(n2650),  .B(n5986),  .C(n5987), .Y(k_data[20]));
   AOI22X1 U7150 ( .A(n2716),  .B(n2955),  .C(n5934),  .D(n2893), .Y(n5989));
   AOI22X1 U7151 ( .A(n5846),  .B(n2956),  .C(n5925),  .D(n5763), .Y(n5988));
   NOR3X1 U7152 ( .A(n2534),  .B(n5853),  .C(n5991), .Y(n5986));
   AOI21X1 U7153 ( .A(n2953),  .B(n2843),  .C(n5899), .Y(n5990));
   AOI22X1 U7154 ( .A(n6001),  .B(n5992),  .C(n5917),  .D(n5993), .Y(n5985));
   OAI21X1 U7155 ( .A(n5899),  .B(n2888),  .C(n5999), .Y(n5997));
   OAI21X1 U7156 ( .A(n5875),  .B(n5993),  .C(n5917), .Y(n5999));
   OAI21X1 U7157 ( .A(n4705),  .B(n2594),  .C(n2782), .Y(n5993));
   NAND3X1 U7158 ( .A(n2845),  .B(n2653),  .C(n1968), .Y(n5996));
   AOI22X1 U7159 ( .A(n5789),  .B(n5885),  .C(n5807),  .D(n5763), .Y(n5995));
   AOI21X1 U7160 ( .A(n5886),  .B(n6021),  .C(n5774), .Y(n5994));
   OAI21X1 U7161 ( .A(n2849),  .B(n2718),  .C(n6004), .Y(n5774));
   AOI22X1 U7162 ( .A(n5782),  .B(n2784),  .C(n6109),  .D(n6001), .Y(n6004));
   OR2X1 U7163 ( .A(n6005),  .B(n6006), .Y(k_data[19]));
   NAND3X1 U7164 ( .A(n6007),  .B(n6008),  .C(n1927), .Y(n6006));
   AOI21X1 U7165 ( .A(n5845),  .B(n2956),  .C(n1758), .Y(n6009));
   NAND2X1 U7166 ( .A(n5814),  .B(n5917), .Y(n6008));
   AOI22X1 U7167 ( .A(n6109),  .B(n2893),  .C(n5846),  .D(n6001), .Y(n6007));
   NAND3X1 U7168 ( .A(n6010),  .B(n6011),  .C(n1924), .Y(n6005));
   AOI22X1 U7169 ( .A(n5789),  .B(n6013),  .C(n5807),  .D(n2719), .Y(n6012));
   NAND3X1 U7170 ( .A(n2654),  .B(n2116),  .C(n1933), .Y(n6013));
   OAI21X1 U7171 ( .A(n5771),  .B(n2717),  .C(n5763), .Y(n6011));
   AOI21X1 U7172 ( .A(n5925),  .B(t_ctr_reg[5]),  .C(n6089), .Y(n6010));
   NOR3X1 U7173 ( .A(n1939),  .B(n1946),  .C(n1949), .Y(n6017));
   AOI21X1 U7174 ( .A(n5849),  .B(n2715),  .C(n2849), .Y(n6020));
   AOI21X1 U7175 ( .A(n2593),  .B(n2783),  .C(n2657), .Y(n6019));
   NAND3X1 U7176 ( .A(n6022),  .B(n2104),  .C(n6023), .Y(n6018));
   OAI21X1 U7177 ( .A(n5843),  .B(n1970),  .C(n5763), .Y(n6023));
   NAND3X1 U7178 ( .A(n2956),  .B(n4705),  .C(n6000), .Y(n6022));
   AOI21X1 U7179 ( .A(n5782),  .B(n2893),  .C(n6025), .Y(n6016));
   OAI21X1 U7180 ( .A(n5916),  .B(n2953),  .C(n6026), .Y(n6025));
   NAND2X1 U7181 ( .A(n5889),  .B(n5917), .Y(n6026));
   AOI21X1 U7182 ( .A(n5821),  .B(n2955),  .C(n5868), .Y(n6015));
   OAI21X1 U7183 ( .A(n2891),  .B(n2954),  .C(n6027), .Y(n5868));
   NAND2X1 U7184 ( .A(n5914),  .B(n5763), .Y(n6027));
   OR2X1 U7185 ( .A(n6028),  .B(n6029), .Y(k_data[17]));
   NAND3X1 U7186 ( .A(n6030),  .B(n6031),  .C(n1925), .Y(n6029));
   AOI22X1 U7187 ( .A(n5845),  .B(n2656),  .C(n5821),  .D(n5763), .Y(n6032));
   NAND2X1 U7188 ( .A(n5843),  .B(n6001), .Y(n6031));
   AOI22X1 U7189 ( .A(n6068),  .B(n4705),  .C(n5873),  .D(n5874), .Y(n6030));
   NAND3X1 U7190 ( .A(n6033),  .B(n6034),  .C(n1926), .Y(n6028));
   AOI22X1 U7191 ( .A(n5917),  .B(n6036),  .C(n5789),  .D(n6037), .Y(n6035));
   NAND3X1 U7192 ( .A(n2715),  .B(n2889),  .C(n2594), .Y(n6037));
   NAND3X1 U7193 ( .A(n2651),  .B(n2107),  .C(n1934), .Y(n6036));
   OAI21X1 U7194 ( .A(n5788),  .B(n5782),  .C(n2955), .Y(n6034));
   NOR3X1 U7195 ( .A(n6043),  .B(n5981),  .C(n1950), .Y(n6042));
   AOI21X1 U7196 ( .A(n2892),  .B(n2783),  .C(n5916), .Y(n6044));
   OAI21X1 U7197 ( .A(n4703),  .B(n2952),  .C(n6046), .Y(n6043));
   OAI21X1 U7198 ( .A(n5769),  .B(n6109),  .C(n5789), .Y(n6046));
   AOI22X1 U7199 ( .A(n5763),  .B(n6047),  .C(n6001),  .D(n6048), .Y(n6041));
   NAND3X1 U7200 ( .A(n2113),  .B(n2890),  .C(n2844), .Y(n6048));
   NAND3X1 U7201 ( .A(n2107),  .B(n2718),  .C(n5792), .Y(n6047));
   AOI21X1 U7202 ( .A(n5904),  .B(n2784),  .C(n1976), .Y(n6040));
   NAND3X1 U7203 ( .A(n6049),  .B(n2109),  .C(n5898), .Y(n5812));
   INVX1 U7204 ( .A(n5980), .Y(n5898));
   OAI21X1 U7205 ( .A(n4705),  .B(n1964),  .C(n2111), .Y(n5980));
   NAND2X1 U7206 ( .A(n5934),  .B(n5886), .Y(n6049));
   NAND3X1 U7207 ( .A(n6051),  .B(n6052),  .C(n6053), .Y(k_data[15]));
   AND2X1 U7208 ( .A(n6054),  .B(n6055), .Y(n6053));
   AOI21X1 U7209 ( .A(n2956),  .B(n5782),  .C(n5959), .Y(n6055));
   OAI21X1 U7210 ( .A(n2847),  .B(n2891),  .C(n6056), .Y(n5959));
   AOI22X1 U7211 ( .A(n5873),  .B(n5874),  .C(n5821),  .D(n2785), .Y(n6056));
   INVX1 U7212 ( .A(n6057), .Y(n6054));
   OAI21X1 U7213 ( .A(n5816),  .B(n2954),  .C(n6058), .Y(n6057));
   AOI22X1 U7214 ( .A(n5934),  .B(n5886),  .C(n5763),  .D(n2846), .Y(n6058));
   NOR3X1 U7215 ( .A(n1940),  .B(n6050),  .C(n6045), .Y(n6052));
   AOI21X1 U7216 ( .A(n5848),  .B(n2103),  .C(n2116), .Y(n6059));
   AOI22X1 U7217 ( .A(n5789),  .B(n6060),  .C(n5772),  .D(n2719), .Y(n6051));
   OAI21X1 U7218 ( .A(n4703),  .B(n2536),  .C(n2889), .Y(n6060));
   OAI21X1 U7219 ( .A(n5861),  .B(n5949),  .C(n6066), .Y(n6065));
   OAI21X1 U7220 ( .A(n5821),  .B(n5767),  .C(n5917), .Y(n6066));
   OAI21X1 U7221 ( .A(n4707),  .B(n2890),  .C(n2842), .Y(n5767));
   NAND3X1 U7222 ( .A(n1955),  .B(n2105),  .C(n1967), .Y(n6064));
   AOI22X1 U7223 ( .A(n5789),  .B(n6070),  .C(n5763),  .D(n2110), .Y(n6063));
   INVX1 U7224 ( .A(n1956), .Y(n6070));
   AOI21X1 U7225 ( .A(n5772),  .B(n6001),  .C(n1851), .Y(n6062));
   AOI22X1 U7226 ( .A(n5934),  .B(n5917),  .C(n5845),  .D(n5789), .Y(n6073));
   AOI22X1 U7227 ( .A(n6050),  .B(n4705),  .C(n5886),  .D(n2591), .Y(n6072));
   AOI21X1 U7228 ( .A(n5789),  .B(n1977),  .C(n5991), .Y(n6079));
   AOI22X1 U7229 ( .A(n5769),  .B(n2719),  .C(n5845),  .D(n2656), .Y(n6078));
   AOI22X1 U7230 ( .A(n5860),  .B(n5917),  .C(n5763),  .D(n2716), .Y(n6076));
   AOI21X1 U7231 ( .A(n5771),  .B(n6001),  .C(n1954), .Y(n6075));
   NAND3X1 U7232 ( .A(n1971),  .B(n2105),  .C(n1928), .Y(n5801));
   AOI21X1 U7233 ( .A(n5807),  .B(n5763),  .C(n1758), .Y(n6081));
   AOI21X1 U7234 ( .A(n5789),  .B(n5992),  .C(n6084), .Y(n6083));
   OAI21X1 U7235 ( .A(n5971),  .B(n2891),  .C(n2712), .Y(n6084));
   OAI21X1 U7236 ( .A(n2782),  .B(n4705),  .C(n2847), .Y(n5992));
   MUX2X1 U7237 ( .A(n5813),  .B(n5886),  .S(n4705), .Y(n6082));
   INVX1 U7238 ( .A(n1961), .Y(n5813));
   AOI21X1 U7239 ( .A(n5917),  .B(n6109),  .C(n6068), .Y(n5865));
   INVX1 U7240 ( .A(n6085), .Y(k_data[12]));
   NOR3X1 U7241 ( .A(n1853),  .B(n1947),  .C(n1951), .Y(n6085));
   NAND3X1 U7242 ( .A(n1971),  .B(n2112),  .C(n6088), .Y(n6087));
   OAI21X1 U7243 ( .A(n5918),  .B(n5771),  .C(n5789), .Y(n6088));
   NAND3X1 U7244 ( .A(n2479),  .B(n2778),  .C(n2845), .Y(n6086));
   NAND3X1 U7245 ( .A(n5763),  .B(t_ctr_reg[3]),  .C(n5859), .Y(n5963));
   AOI22X1 U7246 ( .A(n5917),  .B(n5867),  .C(n5821),  .D(n2956), .Y(n6091));
   AOI22X1 U7247 ( .A(n5783),  .B(t_ctr_reg[3]),  .C(n5873),  .D(n6021), .Y(n6090));
   AND2X1 U7248 ( .A(n6001),  .B(n4707), .Y(n5873));
   NAND3X1 U7249 ( .A(n6092),  .B(n6093),  .C(n6094), .Y(k_data[11]));
   AOI21X1 U7250 ( .A(n2956),  .B(n5934),  .C(n5945), .Y(n6096));
   OAI21X1 U7251 ( .A(n2849),  .B(n2890),  .C(n6097), .Y(n5945));
   AOI22X1 U7252 ( .A(n6069),  .B(n5859),  .C(n5846),  .D(n6001), .Y(n6097));
   INVX1 U7253 ( .A(n6098), .Y(n6095));
   OAI21X1 U7254 ( .A(n5916),  .B(n2892),  .C(n6099), .Y(n6098));
   AOI22X1 U7255 ( .A(n5886),  .B(n6021),  .C(n5771),  .D(n2848), .Y(n6099));
   NOR3X1 U7256 ( .A(n5880),  .B(n5803),  .C(n5991), .Y(n6093));
   AND2X1 U7257 ( .A(n5925),  .B(n5917), .Y(n5880));
   AOI21X1 U7258 ( .A(n5807),  .B(n5917),  .C(n6100), .Y(n6092));
   OAI21X1 U7259 ( .A(n5816),  .B(n2888),  .C(n6101), .Y(n6100));
   OAI21X1 U7260 ( .A(n5788),  .B(n5845),  .C(n5789), .Y(n6101));
   AOI22X1 U7261 ( .A(n5781),  .B(t_ctr_reg[3]),  .C(n5789),  .D(n2108), .Y(n6106));
   AOI22X1 U7262 ( .A(n5821),  .B(n2848),  .C(n2784),  .D(n2717), .Y(n6105));
   NOR3X1 U7263 ( .A(n1943),  .B(n6089),  .C(n1952), .Y(n6103));
   AOI21X1 U7264 ( .A(n2115),  .B(n2106),  .C(n5786), .Y(n6108));
   AOI21X1 U7265 ( .A(n1956),  .B(n2114),  .C(n2720), .Y(n6107));
   AOI21X1 U7266 ( .A(n2716),  .B(t_ctr_reg[3]),  .C(n5918), .Y(n6071));
   AOI22X1 U7267 ( .A(n6001),  .B(n6110),  .C(n5972),  .D(n2955), .Y(n6102));
   OAI21X1 U7268 ( .A(t_ctr_reg[3]),  .B(n5915),  .C(n2847), .Y(n6110));
   OR2X1 U7269 ( .A(n6111),  .B(n6112), .Y(k_data[0]));
   NAND3X1 U7270 ( .A(n6113),  .B(n6114),  .C(n1929), .Y(n6112));
   AOI21X1 U7271 ( .A(n5821),  .B(n6001),  .C(n5953), .Y(n6115));
   OAI21X1 U7272 ( .A(n2849),  .B(n2116),  .C(n6116), .Y(n5953));
   AOI21X1 U7273 ( .A(n5788),  .B(n6001),  .C(n6003), .Y(n6116));
   NAND2X1 U7274 ( .A(n6061),  .B(n2893), .Y(n6114));
   AOI22X1 U7275 ( .A(n5886),  .B(n5885),  .C(n5845),  .D(n2719), .Y(n6113));
   NAND3X1 U7276 ( .A(n6119),  .B(n6120),  .C(n6121), .Y(n6111));
   NOR3X1 U7277 ( .A(n1944),  .B(n6050),  .C(n5912), .Y(n6121));
   NOR3X1 U7278 ( .A(n4703),  .B(t_ctr_reg[4]),  .C(n4711), .Y(n6118));
   AOI21X1 U7279 ( .A(n5832),  .B(n2892),  .C(n2849), .Y(n6122));
   NOR3X1 U7280 ( .A(t_ctr_reg[2]),  .B(t_ctr_reg[3]),  .C(n4707), .Y(n6117));
   AND2X1 U7281 ( .A(n2098),  .B(n2113), .Y(n5832));
   NAND2X1 U7282 ( .A(n5917),  .B(n1970), .Y(n6120));
   INVX1 U7283 ( .A(t_ctr_reg[4]), .Y(n4707));
   AND2X1 U7284 ( .A(t_ctr_reg[2]),  .B(n4711), .Y(n5805));
   INVX1 U7285 ( .A(t_ctr_reg[5]), .Y(n4711));
   INVX1 U7286 ( .A(t_ctr_reg[0]), .Y(n4700));
   AOI22X1 U7287 ( .A(n6068),  .B(n4705),  .C(n5763),  .D(n1979), .Y(n6119));
   INVX1 U7288 ( .A(t_ctr_reg[2]), .Y(n4703));
   INVX1 U7289 ( .A(t_ctr_reg[1]), .Y(n4701));
   INVX1 U7290 ( .A(t_ctr_reg[3]), .Y(n4705));
   OAI21X1 U7291 ( .A(n6123),  .B(n5544),  .C(n6124), .Y(N999));
   OAI21X1 U7292 ( .A(a_reg[30]),  .B(b_reg[30]),  .C(c_reg[30]), .Y(n6124));
   INVX1 U7293 ( .A(b_reg[30]), .Y(n5544));
   OAI21X1 U7294 ( .A(n5418),  .B(n6125),  .C(n6126), .Y(N998));
   OAI21X1 U7295 ( .A(a_reg[31]),  .B(b_reg[31]),  .C(c_reg[31]), .Y(n6126));
   INVX1 U7296 ( .A(b_reg[31]), .Y(n6125));
   FAX1 U7297 ( .A(n4672),  .B(n5400),  .C(a_reg[13]), .YS(N997));
   FAX1 U7298 ( .A(n5362),  .B(n5402),  .C(a_reg[14]), .YS(N996));
   FAX1 U7299 ( .A(n5364),  .B(n5404),  .C(a_reg[15]), .YS(N995));
   FAX1 U7300 ( .A(n6127),  .B(n4681),  .C(a_reg[16]), .YS(N994));
   FAX1 U7301 ( .A(n6128),  .B(n5408),  .C(a_reg[17]), .YS(N993));
   FAX1 U7302 ( .A(n5370),  .B(n4684),  .C(a_reg[18]), .YS(N992));
   FAX1 U7303 ( .A(n5372),  .B(n5412),  .C(a_reg[19]), .YS(N991));
   FAX1 U7304 ( .A(n4675),  .B(n4687),  .C(a_reg[20]), .YS(N990));
   FAX1 U7305 ( .A(n6123),  .B(n5398),  .C(a_reg[10]), .YS(N989));
   FAX1 U7306 ( .A(n5418),  .B(n5400),  .C(a_reg[11]), .YS(N988));
   FAX1 U7307 ( .A(n5402),  .B(n5380),  .C(a_reg[0]), .YS(N987));
   FAX1 U7308 ( .A(n5404),  .B(n6129),  .C(a_reg[13]), .YS(N986));
   FAX1 U7309 ( .A(n4672),  .B(n4681),  .C(a_reg[14]), .YS(N985));
   FAX1 U7310 ( .A(n5362),  .B(n5408),  .C(a_reg[15]), .YS(N984));
   FAX1 U7311 ( .A(n5364),  .B(n4684),  .C(a_reg[16]), .YS(N983));
   FAX1 U7312 ( .A(n6127),  .B(n5412),  .C(a_reg[17]), .YS(N982));
   FAX1 U7313 ( .A(n6128),  .B(n4687),  .C(a_reg[18]), .YS(N981));
   FAX1 U7314 ( .A(n5370),  .B(n6123),  .C(a_reg[19]), .YS(N980));
   FAX1 U7315 ( .A(n5372),  .B(n5418),  .C(a_reg[20]), .YS(N979));
   FAX1 U7316 ( .A(n4675),  .B(n5398),  .C(a_reg[0]), .YS(N978));
   FAX1 U7317 ( .A(n5400),  .B(n6129),  .C(a_reg[10]), .YS(N977));
   FAX1 U7318 ( .A(n4672),  .B(n5402),  .C(a_reg[11]), .YS(N976));
   INVX1 U7319 ( .A(a_reg[2]), .Y(n4672));
   FAX1 U7320 ( .A(n5362),  .B(n5404),  .C(a_reg[12]), .YS(N975));
   FAX1 U7321 ( .A(n5364),  .B(n4681),  .C(a_reg[13]), .YS(N974));
   INVX1 U7322 ( .A(a_reg[25]), .Y(n4681));
   FAX1 U7323 ( .A(n6127),  .B(n5408),  .C(a_reg[14]), .YS(N973));
   FAX1 U7324 ( .A(n6128),  .B(n4684),  .C(a_reg[15]), .YS(N972));
   INVX1 U7325 ( .A(a_reg[27]), .Y(n4684));
   FAX1 U7326 ( .A(n5370),  .B(n5412),  .C(a_reg[16]), .YS(N971));
   FAX1 U7327 ( .A(n5372),  .B(n4687),  .C(a_reg[17]), .YS(N970));
   INVX1 U7328 ( .A(a_reg[29]), .Y(n4687));
   FAX1 U7329 ( .A(n4675),  .B(n6123),  .C(a_reg[18]), .YS(N969));
   INVX1 U7330 ( .A(a_reg[30]), .Y(n6123));
   INVX1 U7331 ( .A(a_reg[9]), .Y(n4675));
   FAX1 U7332 ( .A(n5418),  .B(n6130),  .C(a_reg[10]), .YS(N968));
   INVX1 U7333 ( .A(a_reg[31]), .Y(n5418));
   FAX1 U7334 ( .A(n5396),  .B(n5378),  .C(a_reg[0]), .YS(N967));
   FAX1 U7335 ( .A(n5398),  .B(n6129),  .C(a_reg[12]), .YS(N966));
   INVX1 U7336 ( .A(n6131), .Y(N869));
   MUX2X1 U7337 ( .A(f_reg[0]),  .B(g_reg[0]),  .S(e_reg[0]), .Y(n6131));
   INVX1 U7338 ( .A(n6132), .Y(N868));
   MUX2X1 U7339 ( .A(f_reg[1]),  .B(g_reg[1]),  .S(e_reg[1]), .Y(n6132));
   INVX1 U7340 ( .A(n6133), .Y(N867));
   MUX2X1 U7341 ( .A(f_reg[2]),  .B(g_reg[2]),  .S(e_reg[2]), .Y(n6133));
   INVX1 U7342 ( .A(n6134), .Y(N866));
   MUX2X1 U7343 ( .A(f_reg[3]),  .B(g_reg[3]),  .S(e_reg[3]), .Y(n6134));
   MUX2X1 U7344 ( .A(n4980),  .B(n5108),  .S(e_reg[4]), .Y(N865));
   INVX1 U7345 ( .A(f_reg[4]), .Y(n4980));
   INVX1 U7346 ( .A(g_reg[4]), .Y(n5108));
   INVX1 U7347 ( .A(n6135), .Y(N864));
   MUX2X1 U7348 ( .A(f_reg[5]),  .B(g_reg[5]),  .S(e_reg[5]), .Y(n6135));
   MUX2X1 U7349 ( .A(n4984),  .B(n5112),  .S(e_reg[6]), .Y(N863));
   INVX1 U7350 ( .A(f_reg[6]), .Y(n4984));
   INVX1 U7351 ( .A(g_reg[6]), .Y(n5112));
   INVX1 U7352 ( .A(n6136), .Y(N862));
   MUX2X1 U7353 ( .A(g_reg[7]),  .B(f_reg[7]),  .S(n4858), .Y(n6136));
   INVX1 U7354 ( .A(n6137), .Y(N861));
   MUX2X1 U7355 ( .A(g_reg[8]),  .B(f_reg[8]),  .S(n4860), .Y(n6137));
   MUX2X1 U7356 ( .A(n4990),  .B(n5118),  .S(e_reg[9]), .Y(N860));
   INVX1 U7357 ( .A(f_reg[9]), .Y(n4990));
   INVX1 U7358 ( .A(g_reg[9]), .Y(n5118));
   MUX2X1 U7359 ( .A(n5120),  .B(n4992),  .S(n4864), .Y(N859));
   INVX1 U7360 ( .A(g_reg[10]), .Y(n5120));
   INVX1 U7361 ( .A(f_reg[10]), .Y(n4992));
   INVX1 U7362 ( .A(n6138), .Y(N858));
   MUX2X1 U7363 ( .A(g_reg[11]),  .B(f_reg[11]),  .S(n4866), .Y(n6138));
   INVX1 U7364 ( .A(n6139), .Y(N857));
   MUX2X1 U7365 ( .A(f_reg[12]),  .B(g_reg[12]),  .S(e_reg[12]), .Y(n6139));
   INVX1 U7366 ( .A(n6140), .Y(N856));
   MUX2X1 U7367 ( .A(g_reg[13]),  .B(f_reg[13]),  .S(n4870), .Y(n6140));
   INVX1 U7368 ( .A(e_reg[13]), .Y(n4870));
   INVX1 U7369 ( .A(n6141), .Y(N855));
   MUX2X1 U7370 ( .A(f_reg[14]),  .B(g_reg[14]),  .S(e_reg[14]), .Y(n6141));
   INVX1 U7371 ( .A(n6142), .Y(N854));
   MUX2X1 U7372 ( .A(g_reg[15]),  .B(f_reg[15]),  .S(n4874), .Y(n6142));
   INVX1 U7373 ( .A(n6143), .Y(N853));
   MUX2X1 U7374 ( .A(g_reg[16]),  .B(f_reg[16]),  .S(n4876), .Y(n6143));
   INVX1 U7375 ( .A(n6144), .Y(N852));
   MUX2X1 U7376 ( .A(f_reg[17]),  .B(g_reg[17]),  .S(e_reg[17]), .Y(n6144));
   INVX1 U7377 ( .A(n6145), .Y(N851));
   MUX2X1 U7378 ( .A(f_reg[18]),  .B(g_reg[18]),  .S(e_reg[18]), .Y(n6145));
   MUX2X1 U7379 ( .A(n5010),  .B(n5138),  .S(e_reg[19]), .Y(N850));
   INVX1 U7380 ( .A(f_reg[19]), .Y(n5010));
   INVX1 U7381 ( .A(g_reg[19]), .Y(n5138));
   MUX2X1 U7382 ( .A(n5140),  .B(n5012),  .S(n4884), .Y(N849));
   INVX1 U7383 ( .A(g_reg[20]), .Y(n5140));
   INVX1 U7384 ( .A(f_reg[20]), .Y(n5012));
   MUX2X1 U7385 ( .A(n5142),  .B(n5014),  .S(n4886), .Y(N848));
   INVX1 U7386 ( .A(g_reg[21]), .Y(n5142));
   INVX1 U7387 ( .A(f_reg[21]), .Y(n5014));
   MUX2X1 U7388 ( .A(n5144),  .B(n5016),  .S(n4888), .Y(N847));
   INVX1 U7389 ( .A(g_reg[22]), .Y(n5144));
   INVX1 U7390 ( .A(f_reg[22]), .Y(n5016));
   INVX1 U7391 ( .A(n6146), .Y(N846));
   MUX2X1 U7392 ( .A(g_reg[23]),  .B(f_reg[23]),  .S(n4890), .Y(n6146));
   INVX1 U7393 ( .A(n6147), .Y(N845));
   MUX2X1 U7394 ( .A(f_reg[24]),  .B(g_reg[24]),  .S(e_reg[24]), .Y(n6147));
   INVX1 U7395 ( .A(n6148), .Y(N844));
   MUX2X1 U7396 ( .A(g_reg[25]),  .B(f_reg[25]),  .S(n4894), .Y(n6148));
   INVX1 U7397 ( .A(n6149), .Y(N843));
   MUX2X1 U7398 ( .A(g_reg[26]),  .B(f_reg[26]),  .S(n4896), .Y(n6149));
   INVX1 U7399 ( .A(n6150), .Y(N842));
   MUX2X1 U7400 ( .A(g_reg[27]),  .B(f_reg[27]),  .S(n4898), .Y(n6150));
   INVX1 U7401 ( .A(n6151), .Y(N841));
   MUX2X1 U7402 ( .A(f_reg[28]),  .B(g_reg[28]),  .S(e_reg[28]), .Y(n6151));
   MUX2X1 U7403 ( .A(n5158),  .B(n5030),  .S(n4902), .Y(N840));
   INVX1 U7404 ( .A(g_reg[29]), .Y(n5158));
   INVX1 U7405 ( .A(f_reg[29]), .Y(n5030));
   MUX2X1 U7406 ( .A(n5032),  .B(n5160),  .S(e_reg[30]), .Y(N839));
   INVX1 U7407 ( .A(f_reg[30]), .Y(n5032));
   INVX1 U7408 ( .A(g_reg[30]), .Y(n5160));
   INVX1 U7409 ( .A(n6152), .Y(N838));
   MUX2X1 U7410 ( .A(g_reg[31]),  .B(f_reg[31]),  .S(n4906), .Y(n6152));
   FAX1 U7411 ( .A(e_reg[6]),  .B(n4894),  .C(n4866), .YS(N837));
   FAX1 U7412 ( .A(n4858),  .B(n4896),  .C(e_reg[12]), .YS(N836));
   FAX1 U7413 ( .A(n4860),  .B(n4898),  .C(e_reg[13]), .YS(N835));
   FAX1 U7414 ( .A(e_reg[9]),  .B(e_reg[28]),  .C(e_reg[14]), .YS(N834));
   FAX1 U7415 ( .A(n4902),  .B(n4874),  .C(e_reg[10]), .YS(N833));
   FAX1 U7416 ( .A(e_reg[30]),  .B(n4876),  .C(n4866), .YS(N832));
   FAX1 U7417 ( .A(e_reg[31]),  .B(e_reg[17]),  .C(e_reg[12]), .YS(N831));
   FAX1 U7418 ( .A(e_reg[18]),  .B(e_reg[13]),  .C(e_reg[0]), .YS(N830));
   FAX1 U7419 ( .A(e_reg[1]),  .B(e_reg[19]),  .C(e_reg[14]), .YS(N829));
   FAX1 U7420 ( .A(e_reg[2]),  .B(n4884),  .C(n4874), .YS(N828));
   INVX1 U7421 ( .A(e_reg[15]), .Y(n4874));
   INVX1 U7422 ( .A(e_reg[20]), .Y(n4884));
   FAX1 U7423 ( .A(e_reg[3]),  .B(n4886),  .C(n4876), .YS(N827));
   FAX1 U7424 ( .A(e_reg[4]),  .B(e_reg[22]),  .C(e_reg[17]), .YS(N826));
   FAX1 U7425 ( .A(e_reg[5]),  .B(e_reg[23]),  .C(e_reg[18]), .YS(N825));
   FAX1 U7426 ( .A(e_reg[6]),  .B(e_reg[24]),  .C(e_reg[19]), .YS(N824));
   FAX1 U7427 ( .A(n4858),  .B(n4894),  .C(e_reg[20]), .YS(N823));
   INVX1 U7428 ( .A(e_reg[25]), .Y(n4894));
   FAX1 U7429 ( .A(n4860),  .B(n4896),  .C(e_reg[21]), .YS(N822));
   FAX1 U7430 ( .A(e_reg[9]),  .B(n4898),  .C(n4888), .YS(N821));
   INVX1 U7431 ( .A(e_reg[27]), .Y(n4898));
   FAX1 U7432 ( .A(e_reg[28]),  .B(n4890),  .C(n4864), .YS(N820));
   INVX1 U7433 ( .A(e_reg[10]), .Y(n4864));
   INVX1 U7434 ( .A(e_reg[23]), .Y(n4890));
   FAX1 U7435 ( .A(n4902),  .B(e_reg[24]),  .C(n4866), .YS(N819));
   INVX1 U7436 ( .A(e_reg[11]), .Y(n4866));
   FAX1 U7437 ( .A(e_reg[30]),  .B(e_reg[25]),  .C(e_reg[12]), .YS(N818));
   FAX1 U7438 ( .A(n4906),  .B(n4896),  .C(e_reg[13]), .YS(N817));
   INVX1 U7439 ( .A(e_reg[26]), .Y(n4896));
   INVX1 U7440 ( .A(e_reg[31]), .Y(n4906));
   FAX1 U7441 ( .A(e_reg[27]),  .B(e_reg[14]),  .C(e_reg[0]), .YS(N816));
   FAX1 U7442 ( .A(e_reg[28]),  .B(e_reg[1]),  .C(e_reg[15]), .YS(N815));
   FAX1 U7443 ( .A(e_reg[2]),  .B(n4902),  .C(n4876), .YS(N814));
   INVX1 U7444 ( .A(e_reg[16]), .Y(n4876));
   INVX1 U7445 ( .A(e_reg[29]), .Y(n4902));
   FAX1 U7446 ( .A(e_reg[3]),  .B(e_reg[30]),  .C(e_reg[17]), .YS(N813));
   FAX1 U7447 ( .A(e_reg[4]),  .B(e_reg[31]),  .C(e_reg[18]), .YS(N812));
   FAX1 U7448 ( .A(e_reg[5]),  .B(e_reg[19]),  .C(e_reg[0]), .YS(N811));
   FAX1 U7449 ( .A(e_reg[6]),  .B(e_reg[20]),  .C(e_reg[1]), .YS(N810));
   FAX1 U7450 ( .A(n4858),  .B(e_reg[2]),  .C(n4886), .YS(N809));
   INVX1 U7451 ( .A(e_reg[21]), .Y(n4886));
   INVX1 U7452 ( .A(e_reg[7]), .Y(n4858));
   FAX1 U7453 ( .A(n4860),  .B(e_reg[3]),  .C(n4888), .YS(N808));
   INVX1 U7454 ( .A(e_reg[22]), .Y(n4888));
   INVX1 U7455 ( .A(e_reg[8]), .Y(n4860));
   FAX1 U7456 ( .A(e_reg[9]),  .B(e_reg[4]),  .C(e_reg[23]), .YS(N807));
   FAX1 U7457 ( .A(e_reg[5]),  .B(e_reg[24]),  .C(e_reg[10]), .YS(N806));
   OAI21X1 U7458 ( .A(n6153),  .B(n6154),  .C(n6155), .Y(N1029));
   OAI21X1 U7459 ( .A(a_reg[0]),  .B(b_reg[0]),  .C(c_reg[0]), .Y(n6155));
   INVX1 U7460 ( .A(b_reg[0]), .Y(n6154));
   INVX1 U7461 ( .A(a_reg[0]), .Y(n6153));
   OAI21X1 U7462 ( .A(n6129),  .B(n5486),  .C(n6156), .Y(N1028));
   OAI21X1 U7463 ( .A(a_reg[1]),  .B(b_reg[1]),  .C(c_reg[1]), .Y(n6156));
   INVX1 U7464 ( .A(b_reg[1]), .Y(n5486));
   INVX1 U7465 ( .A(a_reg[1]), .Y(n6129));
   OAI21X1 U7466 ( .A(n5362),  .B(n5490),  .C(n6157), .Y(N1026));
   OAI21X1 U7467 ( .A(a_reg[3]),  .B(b_reg[3]),  .C(c_reg[3]), .Y(n6157));
   INVX1 U7468 ( .A(b_reg[3]), .Y(n5490));
   INVX1 U7469 ( .A(a_reg[3]), .Y(n5362));
   OAI21X1 U7470 ( .A(n5364),  .B(n5492),  .C(n6158), .Y(N1025));
   OAI21X1 U7471 ( .A(a_reg[4]),  .B(b_reg[4]),  .C(c_reg[4]), .Y(n6158));
   INVX1 U7472 ( .A(b_reg[4]), .Y(n5492));
   INVX1 U7473 ( .A(a_reg[4]), .Y(n5364));
   OAI21X1 U7474 ( .A(n6127),  .B(n5494),  .C(n6159), .Y(N1024));
   OAI21X1 U7475 ( .A(a_reg[5]),  .B(b_reg[5]),  .C(c_reg[5]), .Y(n6159));
   INVX1 U7476 ( .A(b_reg[5]), .Y(n5494));
   INVX1 U7477 ( .A(a_reg[5]), .Y(n6127));
   OAI21X1 U7478 ( .A(n6128),  .B(n5496),  .C(n6160), .Y(puf_15_wire_3));
   OAI21X1 U7479 ( .A(a_reg[6]),  .B(b_reg[6]),  .C(c_reg[6]), .Y(n6160));
   INVX1 U7480 ( .A(b_reg[6]), .Y(n5496));
   INVX1 U7481 ( .A(a_reg[6]), .Y(n6128));
   OAI21X1 U7482 ( .A(n5370),  .B(n6161),  .C(n6162), .Y(N1022));
   OAI21X1 U7483 ( .A(a_reg[7]),  .B(b_reg[7]),  .C(c_reg[7]), .Y(n6162));
   INVX1 U7484 ( .A(b_reg[7]), .Y(n6161));
   INVX1 U7485 ( .A(a_reg[7]), .Y(n5370));
   OAI21X1 U7486 ( .A(n5372),  .B(n5500),  .C(n6163), .Y(N1021));
   OAI21X1 U7487 ( .A(a_reg[8]),  .B(b_reg[8]),  .C(c_reg[8]), .Y(n6163));
   INVX1 U7488 ( .A(b_reg[8]), .Y(n5500));
   INVX1 U7489 ( .A(a_reg[8]), .Y(n5372));
   OAI21X1 U7490 ( .A(n5378),  .B(n6164),  .C(n6165), .Y(N1018));
   OAI21X1 U7491 ( .A(a_reg[11]),  .B(b_reg[11]),  .C(c_reg[11]), .Y(n6165));
   INVX1 U7492 ( .A(b_reg[11]), .Y(n6164));
   INVX1 U7493 ( .A(a_reg[11]), .Y(n5378));
   OAI21X1 U7494 ( .A(n5380),  .B(n5508),  .C(n6166), .Y(N1017));
   OAI21X1 U7495 ( .A(a_reg[12]),  .B(b_reg[12]),  .C(c_reg[12]), .Y(n6166));
   INVX1 U7496 ( .A(b_reg[12]), .Y(n5508));
   INVX1 U7497 ( .A(a_reg[12]), .Y(n5380));
   OAI21X1 U7498 ( .A(n6167),  .B(n6168),  .C(n6169), .Y(N1016));
   OAI21X1 U7499 ( .A(a_reg[13]),  .B(b_reg[13]),  .C(c_reg[13]), .Y(n6169));
   INVX1 U7500 ( .A(b_reg[13]), .Y(n6168));
   INVX1 U7501 ( .A(a_reg[13]), .Y(n6167));
   OAI21X1 U7502 ( .A(n6170),  .B(n5512),  .C(n6171), .Y(N1015));
   OAI21X1 U7503 ( .A(a_reg[14]),  .B(b_reg[14]),  .C(c_reg[14]), .Y(n6171));
   INVX1 U7504 ( .A(b_reg[14]), .Y(n5512));
   INVX1 U7505 ( .A(a_reg[14]), .Y(n6170));
   OAI21X1 U7506 ( .A(n6172),  .B(n6173),  .C(n6174), .Y(N1014));
   OAI21X1 U7507 ( .A(a_reg[15]),  .B(b_reg[15]),  .C(c_reg[15]), .Y(n6174));
   INVX1 U7508 ( .A(b_reg[15]), .Y(n6173));
   INVX1 U7509 ( .A(a_reg[15]), .Y(n6172));
   OAI21X1 U7510 ( .A(n6175),  .B(n6176),  .C(n6177), .Y(N1013));
   OAI21X1 U7511 ( .A(a_reg[16]),  .B(b_reg[16]),  .C(c_reg[16]), .Y(n6177));
   INVX1 U7512 ( .A(b_reg[16]), .Y(n6176));
   INVX1 U7513 ( .A(a_reg[16]), .Y(n6175));
   OAI21X1 U7514 ( .A(n5390),  .B(n6178),  .C(n6179), .Y(N1012));
   OAI21X1 U7515 ( .A(a_reg[17]),  .B(b_reg[17]),  .C(c_reg[17]), .Y(n6179));
   INVX1 U7516 ( .A(b_reg[17]), .Y(n6178));
   INVX1 U7517 ( .A(a_reg[17]), .Y(n5390));
   OAI21X1 U7518 ( .A(n5392),  .B(n6180),  .C(n6181), .Y(N1011));
   OAI21X1 U7519 ( .A(a_reg[18]),  .B(b_reg[18]),  .C(c_reg[18]), .Y(n6181));
   INVX1 U7520 ( .A(b_reg[18]), .Y(n6180));
   INVX1 U7521 ( .A(a_reg[18]), .Y(n5392));
   OAI21X1 U7522 ( .A(n6130),  .B(n5522),  .C(n6182), .Y(N1010));
   OAI21X1 U7523 ( .A(a_reg[19]),  .B(b_reg[19]),  .C(c_reg[19]), .Y(n6182));
   INVX1 U7524 ( .A(b_reg[19]), .Y(n5522));
   INVX1 U7525 ( .A(a_reg[19]), .Y(n6130));
   OAI21X1 U7526 ( .A(n5396),  .B(n5524),  .C(n6183), .Y(N1009));
   OAI21X1 U7527 ( .A(a_reg[20]),  .B(b_reg[20]),  .C(c_reg[20]), .Y(n6183));
   INVX1 U7528 ( .A(b_reg[20]), .Y(n5524));
   INVX1 U7529 ( .A(a_reg[20]), .Y(n5396));
   OAI21X1 U7530 ( .A(n5398),  .B(n6184),  .C(n6185), .Y(N1008));
   OAI21X1 U7531 ( .A(a_reg[21]),  .B(b_reg[21]),  .C(c_reg[21]), .Y(n6185));
   INVX1 U7532 ( .A(b_reg[21]), .Y(n6184));
   INVX1 U7533 ( .A(a_reg[21]), .Y(n5398));
   OAI21X1 U7534 ( .A(n5400),  .B(n6186),  .C(n6187), .Y(N1007));
   OAI21X1 U7535 ( .A(a_reg[22]),  .B(b_reg[22]),  .C(c_reg[22]), .Y(n6187));
   INVX1 U7536 ( .A(b_reg[22]), .Y(n6186));
   INVX1 U7537 ( .A(a_reg[22]), .Y(n5400));
   OAI21X1 U7538 ( .A(n5402),  .B(n5530),  .C(n6188), .Y(N1006));
   OAI21X1 U7539 ( .A(a_reg[23]),  .B(b_reg[23]),  .C(c_reg[23]), .Y(n6188));
   INVX1 U7540 ( .A(b_reg[23]), .Y(n5530));
   INVX1 U7541 ( .A(a_reg[23]), .Y(n5402));
   OAI21X1 U7542 ( .A(n5404),  .B(n6189),  .C(n6190), .Y(N1005));
   OAI21X1 U7543 ( .A(a_reg[24]),  .B(b_reg[24]),  .C(c_reg[24]), .Y(n6190));
   INVX1 U7544 ( .A(b_reg[24]), .Y(n6189));
   INVX1 U7545 ( .A(a_reg[24]), .Y(n5404));
   OAI21X1 U7546 ( .A(n5408),  .B(n5536),  .C(n6191), .Y(N1003));
   OAI21X1 U7547 ( .A(a_reg[26]),  .B(b_reg[26]),  .C(c_reg[26]), .Y(n6191));
   INVX1 U7548 ( .A(b_reg[26]), .Y(n5536));
   INVX1 U7549 ( .A(a_reg[26]), .Y(n5408));
   OAI21X1 U7550 ( .A(n5412),  .B(n6192),  .C(n6193), .Y(N1001));
   OAI21X1 U7551 ( .A(a_reg[28]),  .B(b_reg[28]),  .C(c_reg[28]), .Y(n6193));
   INVX1 U7552 ( .A(b_reg[28]), .Y(n6192));
   INVX1 U7553 ( .A(a_reg[28]), .Y(n5412));
   INVX1 puf_0_instance_0 ( .A(puf_0_wire_1), .Y(puf_0_wire_0));
   INVX1 puf_0_instance_1 ( .A(puf_0_wire_0), .Y(puf_0_wire_1));
   INVX1 puf_0_instance_2 ( .A(puf_0_wire_3), .Y(puf_0_wire_2));
   MUX2X1 puf_0_instance_3 ( .A(puf_0_wire_2),  .B(puf_0_wire_0),  .S(sel), .Y(digest[112]));
   BUFX2 puf_out_instance_0 ( .A(digest[112]), .Y(pufout[0]));
   INVX1 puf_1_instance_0 ( .A(puf_1_wire_1), .Y(puf_1_wire_0));
   INVX1 puf_1_instance_1 ( .A(puf_1_wire_0), .Y(puf_1_wire_1));
   INVX1 puf_1_instance_2 ( .A(puf_1_wire_3), .Y(puf_1_wire_2));
   MUX2X1 puf_1_instance_3 ( .A(puf_1_wire_2),  .B(puf_1_wire_0),  .S(sel), .Y(n1867));
   BUFX2 puf_out_instance_1 ( .A(n1867), .Y(pufout[1]));
   INVX1 puf_2_instance_0 ( .A(puf_2_wire_1), .Y(puf_2_wire_0));
   INVX1 puf_2_instance_1 ( .A(puf_2_wire_0), .Y(puf_2_wire_1));
   INVX1 puf_2_instance_2 ( .A(puf_2_wire_3), .Y(puf_2_wire_2));
   MUX2X1 puf_2_instance_3 ( .A(puf_2_wire_2),  .B(puf_2_wire_0),  .S(sel), .Y(n2006));
   BUFX2 puf_out_instance_2 ( .A(n2006), .Y(pufout[2]));
   INVX1 puf_3_instance_0 ( .A(puf_3_wire_1), .Y(puf_3_wire_0));
   INVX1 puf_3_instance_1 ( .A(puf_3_wire_0), .Y(puf_3_wire_1));
   INVX1 puf_3_instance_2 ( .A(puf_3_wire_3), .Y(puf_3_wire_2));
   MUX2X1 puf_3_instance_3 ( .A(puf_3_wire_2),  .B(puf_3_wire_0),  .S(sel), .Y(n2067));
   BUFX2 puf_out_instance_3 ( .A(n2067), .Y(pufout[3]));
   INVX1 puf_4_instance_0 ( .A(puf_4_wire_1), .Y(puf_4_wire_0));
   INVX1 puf_4_instance_1 ( .A(puf_4_wire_0), .Y(puf_4_wire_1));
   INVX1 puf_4_instance_2 ( .A(puf_4_wire_3), .Y(puf_4_wire_2));
   MUX2X1 puf_4_instance_3 ( .A(puf_4_wire_2),  .B(puf_4_wire_0),  .S(sel), .Y(n2126));
   BUFX2 puf_out_instance_4 ( .A(n2126), .Y(pufout[4]));
   INVX1 puf_5_instance_0 ( .A(puf_5_wire_1), .Y(puf_5_wire_0));
   INVX1 puf_5_instance_1 ( .A(puf_5_wire_0), .Y(puf_5_wire_1));
   INVX1 puf_5_instance_2 ( .A(puf_5_wire_3), .Y(puf_5_wire_2));
   MUX2X1 puf_5_instance_3 ( .A(puf_5_wire_2),  .B(puf_5_wire_0),  .S(sel), .Y(n2287));
   BUFX2 puf_out_instance_5 ( .A(n2287), .Y(pufout[5]));
   INVX1 puf_6_instance_0 ( .A(puf_6_wire_1), .Y(puf_6_wire_0));
   INVX1 puf_6_instance_1 ( .A(puf_6_wire_0), .Y(puf_6_wire_1));
   INVX1 puf_6_instance_2 ( .A(puf_6_wire_3), .Y(puf_6_wire_2));
   MUX2X1 puf_6_instance_3 ( .A(puf_6_wire_2),  .B(puf_6_wire_0),  .S(sel), .Y(n2688));
   BUFX2 puf_out_instance_6 ( .A(n2688), .Y(pufout[6]));
   INVX1 puf_7_instance_0 ( .A(puf_7_wire_1), .Y(puf_7_wire_0));
   INVX1 puf_7_instance_1 ( .A(puf_7_wire_0), .Y(puf_7_wire_1));
   INVX1 puf_7_instance_2 ( .A(puf_7_wire_3), .Y(puf_7_wire_2));
   MUX2X1 puf_7_instance_3 ( .A(puf_7_wire_2),  .B(puf_7_wire_0),  .S(sel), .Y(n2955));
   BUFX2 puf_out_instance_7 ( .A(n2955), .Y(pufout[7]));
   INVX1 puf_8_instance_0 ( .A(puf_8_wire_1), .Y(puf_8_wire_0));
   INVX1 puf_8_instance_1 ( .A(puf_8_wire_0), .Y(puf_8_wire_1));
   INVX1 puf_8_instance_2 ( .A(puf_8_wire_3), .Y(puf_8_wire_2));
   MUX2X1 puf_8_instance_3 ( .A(puf_8_wire_2),  .B(puf_8_wire_0),  .S(sel), .Y(w_mem_inst_n1827));
   BUFX2 puf_out_instance_8 ( .A(w_mem_inst_n1827), .Y(pufout[8]));
   INVX1 puf_9_instance_0 ( .A(puf_9_wire_1), .Y(puf_9_wire_0));
   INVX1 puf_9_instance_1 ( .A(puf_9_wire_0), .Y(puf_9_wire_1));
   INVX1 puf_9_instance_2 ( .A(puf_9_wire_3), .Y(puf_9_wire_2));
   MUX2X1 puf_9_instance_3 ( .A(puf_9_wire_2),  .B(puf_9_wire_0),  .S(sel), .Y(w_mem_inst_n1699));
   BUFX2 puf_out_instance_9 ( .A(w_mem_inst_n1699), .Y(pufout[9]));
   INVX1 puf_10_instance_0 ( .A(puf_10_wire_1), .Y(puf_10_wire_0));
   INVX1 puf_10_instance_1 ( .A(puf_10_wire_0), .Y(puf_10_wire_1));
   INVX1 puf_10_instance_2 ( .A(puf_10_wire_3), .Y(puf_10_wire_2));
   MUX2X1 puf_10_instance_3 ( .A(puf_10_wire_2),  .B(puf_10_wire_0),  .S(sel), .Y(n3445));
   BUFX2 puf_out_instance_10 ( .A(n3445), .Y(pufout[10]));
   INVX1 puf_11_instance_0 ( .A(puf_11_wire_1), .Y(puf_11_wire_0));
   INVX1 puf_11_instance_1 ( .A(puf_11_wire_0), .Y(puf_11_wire_1));
   INVX1 puf_11_instance_2 ( .A(puf_11_wire_3), .Y(puf_11_wire_2));
   MUX2X1 puf_11_instance_3 ( .A(puf_11_wire_2),  .B(puf_11_wire_0),  .S(sel), .Y(n4678));
   BUFX2 puf_out_instance_11 ( .A(n4678), .Y(pufout[11]));
   INVX1 puf_12_instance_0 ( .A(puf_12_wire_1), .Y(puf_12_wire_0));
   INVX1 puf_12_instance_1 ( .A(puf_12_wire_0), .Y(puf_12_wire_1));
   INVX1 puf_12_instance_2 ( .A(puf_12_wire_3), .Y(puf_12_wire_2));
   MUX2X1 puf_12_instance_3 ( .A(puf_12_wire_2),  .B(puf_12_wire_0),  .S(sel), .Y(n1356));
   BUFX2 puf_out_instance_12 ( .A(n1356), .Y(pufout[12]));
   INVX1 puf_13_instance_0 ( .A(puf_13_wire_1), .Y(puf_13_wire_0));
   INVX1 puf_13_instance_1 ( .A(puf_13_wire_0), .Y(puf_13_wire_1));
   INVX1 puf_13_instance_2 ( .A(puf_13_wire_3), .Y(puf_13_wire_2));
   MUX2X1 puf_13_instance_3 ( .A(puf_13_wire_2),  .B(puf_13_wire_0),  .S(sel), .Y(n1336));
   BUFX2 puf_out_instance_13 ( .A(n1336), .Y(pufout[13]));
   INVX1 puf_14_instance_0 ( .A(puf_14_wire_1), .Y(puf_14_wire_0));
   INVX1 puf_14_instance_1 ( .A(puf_14_wire_0), .Y(puf_14_wire_1));
   INVX1 puf_14_instance_2 ( .A(puf_14_wire_3), .Y(puf_14_wire_2));
   MUX2X1 puf_14_instance_3 ( .A(puf_14_wire_2),  .B(puf_14_wire_0),  .S(sel), .Y(n5620));
   BUFX2 puf_out_instance_14 ( .A(n5620), .Y(pufout[14]));
   INVX1 puf_15_instance_0 ( .A(puf_15_wire_1), .Y(puf_15_wire_0));
   INVX1 puf_15_instance_1 ( .A(puf_15_wire_0), .Y(puf_15_wire_1));
   INVX1 puf_15_instance_2 ( .A(puf_15_wire_3), .Y(puf_15_wire_2));
   MUX2X1 puf_15_instance_3 ( .A(puf_15_wire_2),  .B(puf_15_wire_0),  .S(sel), .Y(N1023));
   BUFX2 puf_out_instance_15 ( .A(N1023), .Y(pufout[15]));
endmodule


